/*===========================================*\
Filename         : sgdma_ip.v
Project name     : sgdma_subsys_tst
Description      : Merge all submodules of DMA controller core.
Called by        : sgdma_subsys.v
Email            : bingsong.wang@anlogic.com
Modified         : v1.0 Original version,accomplish the basic functions;20210412	  
Copyright(c)Shanghai Anlu Information Technology Co.,Ltd
\*===========================================*/
`include "../../src/sgdma_ip/def/para_def.vh"
module sgdma_ip(
	input   core_rst_n,
	input   core_clk,
	
	input   [1:0]    lbc_ext_cs_i,
    output  [1:0]    ext_lbc_ack_o,
    input   [31:0]   lbc_ext_addr_i,
    input   [3:0]    lbc_ext_wr_i,
    output  [63:0]   ext_lbc_din_o, 
    input   [31:0]   lbc_ext_dout_i,
	input            lbc_ext_rom_access_i,
	input            lbc_ext_io_access_i,
	input   [2:0]    lbc_ext_bar_num_i,
	input            lbc_ext_vfunc_active_i,
	input   [1:0]    lbc_ext_vfunc_num_i,
	
	output   client0_addr_align_en_o,
	output   [`HEADER_WIDTH-1:0] client0_tlp_header_o,
	output   client0_tlp_dv_o,
	output   client0_tlp_eot_o,
	output   client0_tlp_bad_eot_o,
	output   client0_tlp_hv_o,
	output   [12:0]   client0_tlp_byte_len_o,
	output   [`DATA_WIDTH-1:0]   client0_tlp_data_o,
	output   client0_tlp_func_num_o,
	output   [1:0]   client0_tlp_vfunc_num_o,
	output   client0_tlp_vfunc_active_o,
	input    xadm_client0_halt_i,
	output   client0_tlp_atu_bypass_o,
	
	output   client1_addr_align_en_o,
	output   [`HEADER_WIDTH-1:0] client1_tlp_header_o,
	output   client1_tlp_dv_o,
	output   client1_tlp_eot_o,
	output   client1_tlp_bad_eot_o,
	output   client1_tlp_hv_o,
	output   [12:0]   client1_tlp_byte_len_o,
	output   [`DATA_WIDTH-1:0]   client1_tlp_data_o,
	output   client1_tlp_func_num_o,
	output   [1:0]   client1_tlp_vfunc_num_o,
	output   client1_tlp_vfunc_active_o,
	input    xadm_client1_halt_i,
	output   client1_tlp_atu_bypass_o,
	
	input           radm_bypass_dv_i,
	input           radm_bypass_hv_i,
	input           radm_bypass_eot_i,
	input   [`DATA_WIDTH-1:0]     radm_bypass_data_i,
	input   [`HEADER_WIDTH-1:0]   radm_bypass_header_i,//pos&non_pos 4DW,cpl 3DW. 
	input   [1:0]   radm_bypass_dwen_i,
	input           radm_bypass_cpl_last_i,
	input           radm_bypass_dllp_abort_i,
	input           radm_bypass_tlp_abort_i,
	input           radm_bypass_ecrc_err_i,
	input           radm_bypass_func_num_i,
	input   [1:0]   radm_bypass_vfunc_num_i,
	input           radm_bypass_vfunc_active_i,
	input           radm_bypass_io_req_in_range_i,
	input   [2:0]   radm_bypass_in_membar_range_i,
	input           radm_bypass_rom_in_range_i,
`ifdef AXIL_MBUS0_EN	
	output 	[31:0]   m_axil_awaddr_o,
	output 	[2:0]    m_axil_awprot_o,	
	output 	m_axil_awvalid_o,	
	input  	m_axil_awready_i,	
	output 	[31:0]   m_axil_wdata_o,	
	output 	[3:0]    m_axil_wstrb_o,	
	output 	m_axil_wvalid_o,	
	input  	m_axil_wready_i,	
	input  	m_axil_bvalid_i,	
	input  	[1:0] m_axil_bresp_i,	
	output 	m_axil_bready_o,
	output 	[31:0]   m_axil_araddr_o,	
	output 	[2:0]    m_axil_arprot_o,	
	output 	m_axil_arvalid_o,	
	input  	m_axil_arready_i,	
	input  	[31:0]   m_axil_rdata_i,	
	input  	[1:0]    m_axil_rresp_i,	
	input  	m_axil_rvalid_i,		
	output 	m_axil_rready_o,	
`endif	
`ifdef AXIL_SBUS0_EN
	input   [31:0]   s_axil_awaddr_i,
	input   [2:0]    s_axil_awprot_i,
	input            s_axil_awvalid_i,	
	output           s_axil_awready_o,	
	input   [31:0]   s_axil_wdata_i,	
	input   [3:0]    s_axil_wstrb_i,	
	input            s_axil_wvalid_i,	
	output           s_axil_wready_o,	
	output           s_axil_bvalid_o,	
	output  [1:0]    s_axil_bresp_o,	
	input            s_axil_bready_i,	
	input   [31:0]   s_axil_araddr_i,	
	input   [2:0]    s_axil_arprot_i,	
	input            s_axil_arvalid_i,	
	output           s_axil_arready_o,	
	output  [31:0]   s_axil_rdata_o,	
	output  [1:0]    s_axil_rresp_o,	
	output           s_axil_rvalid_o,	
	input            s_axil_rready_i,
`endif

`ifdef AXIS_BUS0_EN
	output   s0_axis_tx_rst_o,
    output   m0_axis_rx_rst_o,
    output   s0_axis_tx_run_o,
    output   m0_axis_rx_run_o,
    
	output   s0_axis_tx_tready_o,
    input    [`DATA_WIDTH-1:0]    s0_axis_tx_tdata_i,
    input    [`KEEP_WIDTH-1:0]    s0_axis_tx_tkeep_i,
    input    [`KEEP_WIDTH-1:0]    s0_axis_tx_tuser_i,
    input    s0_axis_tx_tlast_i,
    input    s0_axis_tx_tvalid_i,	
	input    m0_axis_rx_tready_i,
    output   [`DATA_WIDTH-1:0]    m0_axis_rx_tdata_o,
    output   [`KEEP_WIDTH-1:0]    m0_axis_rx_tkeep_o,
    output   [`KEEP_WIDTH-1:0]    m0_axis_rx_tuser_o,
    output   m0_axis_rx_tlast_o,
    output   m0_axis_rx_tvalid_o,
`endif
`ifdef AXIS_BUS1_EN
	output   s1_axis_tx_tready_o,
    input    [`DATA_WIDTH-1:0]    s1_axis_tx_tdata_i,
    input    [`KEEP_WIDTH-1:0]    s1_axis_tx_tkeep_i,
    input    [`KEEP_WIDTH-1:0]    s1_axis_tx_tuser_i,
    input    s1_axis_tx_tlast_i,
    input    s1_axis_tx_tvalid_i,
	input    m1_axis_rx_tready_i,
    output   [`DATA_WIDTH-1:0]    m1_axis_rx_tdata_o,
    output   [`KEEP_WIDTH-1:0]    m1_axis_rx_tkeep_o,
    output   [`KEEP_WIDTH-1:0]    m1_axis_rx_tuser_o,
    output   m1_axis_rx_tlast_o,
    output   m1_axis_rx_tvalid_o,
`endif
`ifdef AXI4_BUS0_EN
	input   m_axi_arready_i,
	output  [3:0] m_axi_arid_o,
	output  [`DATA_WIDTH-1:0] m_axi_araddr_o,
	//specifies the number of data transfers that occur within each burst.
	output  [7:0] m_axi_arlen_o,
	//specifies the maximum number of data bytes to transfer in each beat. 011-8byte,100-16byte
	output  [2:0] m_axi_arsize_o,
	output  [1:0] m_axi_arburst_o,
	output  [2:0] m_axi_arprot_o,
	output  m_axi_arvalid_o,
	output  m_axi_arlock_o,
	output  [3:0] m_axi_arcache_o,
	
	input   [3:0] m_axi_rid_i,
	input   [`DATA_WIDTH-1:0]m_axi_rdata_i,
	input   [1:0] m_axi_rresp_i,
	input   m_axi_rlast_i,
	input   m_axi_rvalid_i,
	output  m_axi_rready_o,
	
	input   m_axi_awready_i,
	output  [3:0] m_axi_awid_o,
	output  [`DATA_WIDTH-1:0] m_axi_awaddr_o,
	output  [7:0] m_axi_awlen_o,
	output  [2:0] m_axi_awsize_o,
	output  [1:0] m_axi_awburst_o,
	output  [2:0] m_axi_awprot_o,
	output  m_axi_awvalid_o,
	output  m_axi_awlock_o,
	output  [3:0] m_axi_awcache_o,
	output  [`DATA_WIDTH-1:0] m_axi_wdata_o,
	output  [7:0] m_axi_wstrb_o,
	input   m_axi_wready_i,
	output  m_axi_wlast_o,
	output  m_axi_wvalid_o,
	input   [3:0] m_axi_bid_i,
	input   [1:0] m_axi_bresp_i,
	input   m_axi_bvalid_i,
	output  m_axi_bready_o,
`endif	
`ifdef USR_IRQ_EN
	input   ven_msi_grant_i,
	input   [1:0]   cfg_msi_en_i,
	input   [63:0]  cfg_msi_mask_i,	
	output  ven_msi_req_o,
	output  ven_msi_func_num_o,
	output  [1:0]   ven_msi_vfunc_num_o,
	output  ven_msi_vfunc_active_o,
	output  [2:0]   ven_msi_tc_o,
	output  [4:0]   ven_msi_vector_o,
	output  [63:0]  cfg_msi_pending_o,
	/*
	input   [1:0]    cfg_int_disable_i,
	input   [15:0]   cfg_int_pin_i,
	input   assert_inta_grt_i,
	input   assert_intb_grt_i,
	input   assert_intc_grt_i,
	input   assert_intd_grt_i,
	input   deassert_inta_grt_i,
	input   deassert_intb_grt_i,
	input   deassert_intc_grt_i,
	input   deassert_intd_grt_i,
	output  [1:0]   sys_int_o,
	*/
	input   [`DMA_USR_IRQ-1:0]   usr_irq_req_i,
	output  [`DMA_USR_IRQ-1:0]   usr_irq_ack_o,
	output  msi_enable_o,
	output  [2:0]   msi_vector_width_o,
`endif
//  output                                  rdscp0_eot_out,
//    output                                rd0_rden_out,
`ifdef CFG_MGMT_EN 
	//---dbi2cfg interface---
	input   rdlh_link_up_i,
	output  [31:0]  drp_dbi_din_o,
    output  [3:0]   drp_dbi_wr_o,
    output  [31:0]  drp_dbi_addr_o,
    output 	        drp_dbi_cs_o,
	output          drp_dbi_cs2_o,
    input   [31:0]  drp_lbc_dbi_dout_i,//synthesis keep 
    input 	        drp_lbc_dbi_ack_i, //synthesis keep 
    output  [1:0]   drp_dbi_vfunc_num_o,	
    output          drp_dbi_vfunc_active_o,
	output          drp_dbi_func_num_o,
	output          drp_dbi_rom_access_o,
	output          drp_dbi_io_access_o,
	output          drp_app_dbi_ro_wr_disable_o,
	output  [2:0]   drp_dbi_bar_num_o,	
	input   [18:0]  cfg_mgmt_addr_i,
	input   cfg_mgmt_write_i,
	input   [31:0]  cfg_mgmt_write_data_i,
	input   [3:0]   cfg_mgmt_byte_enable_i,	
	input   cfg_mgmt_read_i,	
	output  [31:0]  cfg_mgmt_read_data_o,	
	output  cfg_mgmt_read_write_done_o,
	input   cfg_mgmt_type1_cfg_reg_access_i
`endif
);
//---Start encrypt;
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-009"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
YBcmXOy/vkPCObchB6FdB+rb39hTDhhwe+0TJLFh2ZbJdUc4ily9fVVeaAkFgNnE
Hpyd4K9wTL2WRsen3ljz78JExJTdpXX2oSjcIofsmb64oX3mUjsIyT1K3TJhznVm
PC3xxPIqHn6ndb/juLRk/OO+TqK9aQaYHnrF313SIgc=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
KemW48uRToqRMyYeirxqg66SEc5eUIB8t6WAuQEDN3S7A+G0IrKr/Vd+SWx5OZ5D
dUv/eNpywhjEDBkyYm8xXcM4iEoCKi5+aOybPmMii7adDJTwLUeQ9n6G6uWHSsX8
jM3OgrsUpP/oj3H6ntu4eNDudozDOtd5EZsfH7wa9ikPlIuogUDcUWI0CMMPA/xY
ei7epFr0t0h90KAdD+ienkAc8pEb+1oN8+KLsbtXZYu8pE1nrMVNxnSJu313Hx3S
u1tWP/9WDrBH5AmaBLzqF4kkBg5AUv+Ekm/mK/p1+ccBPzK26AIO83H++xsVxdqN
Q4Pho1Md3T6fZbxlYT+evw==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
SycmF0xma+RK9LrZqHOR2EK0ajGtoTpm78aPammFf0C1UWJ/H3leNyALKPFaneuP
COklOJDMT5jA+dULOu20QT9XCmp3WXxrNBbs3VQAN8Svji3EO2ECPW68Y7ItfH92
2WKK/LQPwroj6Xb+RxlJhIn5HoiK2Q+PxpAmwQocJ9k=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 353872)
`pragma protect data_block
mCTshtcxo3cJWYEm+3h9GgVAQZHquVMpfY52lnYIYImDLGsS9QV9cvzQQTOKlIKj
8+IIdWhRPgtTbfSnfPrz4tbgBEwB2ezWoi8Sr/XYwg5Ri3/JL5E3lTm2L0GT/dNv
FDp4mAEG7QHwDZ0va+mNdjBNofIlvAy5jWVuxGnSxbzi0/Lt6P2jLVpHNTKJOK13
3uq2Mdz8JHszVooNzj7iFYJAu5Vt631jHODmK2btYoQOrC2nHAwB5K2Nwf7cKMD/
NjqZ9NiS54RL5RpFGEK4Ba5lss4U30yo7377hD+ICR1hukux3cL7BwcYBTBpL6oh
YGPGge8KXVJotn7Y5FeCB0yMhLOb0iOJP/dr/DJ280yVQSyfK0UXtFu1Zdj7aszZ
4S2a8ldIP7Tw9A4VrlOq3ICdFd0zClCIHt/n/U5Axnv/6jtf41q3HvZh90Zl84JT
Et67X6KzXthY/nlWf5iz8DLxKSZu+VaYVHdZFkLiqkz0N0GmZ1zFziNzsljPonQS
eJpgDahLjz61eY8N2U0AAuQbB1/ASkN5gfUYEgxiwC9VAaF+Xb8YCUrRkEciTGjd
SojBw0TUhaO5cKI8HMbXJauylJMJWnH6TDhzay0qQVKrYfLJzbz7ec4ukpXo1veJ
/PW9DZCXiw5dtrBYSNpPhSzpuTyroOWDCLbFOQX3Mwt76+4A85/zgyO0BLJh9x2c
g0quCO6qdvkoZI8f19pV8Lzvi8Xkp32IrAHoBlXSkP0QQ2NqsWkDa843VJxDsd8o
rZDzDKHiRqG27v9t+qftceoKe+TBiG9mfwyOuIq4CNi20c3/DEuLzJ5RZGka2fyz
5S2+oCU/AMY7AuXTLIrJi8L41e0JT76uM+tn65aysP/VTqL6r36TnnSjdcSUgOI7
FMwzLkdvAdUFDNPuULPRXonQSQq42XCuHnKKu70PZ6lCNs/ISKudQgCZyTK4OEQ1
0saucQdbJJq2f84jUYdMW8NS5p33kuVatcJuniZ08x3Te+0XsznPPozXkTSj28IV
k8gToDnqxUxBwvSnS8VvW/lqLeMyRYff2eEGQBhM9cKFYjX7cvJQFS8umpsi/hWq
pFteW1SFwNOqBuR5KTkbiGmOlAqPG8I2mDX77SLDG/fz48fgub8EXOpGKglU5gMU
4rTkeZu0xNa8mcKMrvCmtcqPQVVdVgj+Yf1fPk1d/WDPcRlFVvQgD4Nrjj2ETQwN
69QWyj06KKE7RLuNQpBTumsi+R5CT+2hymrZtNuKHtC/zKprhAd9pCYFU3vbxNj2
aqXHYXhnBrqmzHlucu9DnvM7Q1yEOM6saagsbqtNasNurHTlYEJ78eevtRm7txnr
9xWNHuXzrGbcStAaFV41PBbJvO2b9ZlVOA1M5+/Of6v6nZXiWb6eeaSezf45NRWP
teRSyU+G8yeK4T/nwHqX3iFC2bOe0BvRKQ5z7S8n/BR8iDwy10YAuWmX2l0Szw/u
jQcDRb/UBjkf84/Jcgads+yl5qTvIhrplZ2u6BCA8Bs6RQ+qKro3V55BZVPHkpHo
Df0aEjM3fSuECBNNG6Tv9xgjOz9WHxRYJpXKp4LqiI+uVjMBJJjHlRDCDhbQ/2Dx
MVtzF1LBkadlCYXp/qBYpqi8GItERmonCGXJd8JByhvVkOu8C0srZe6lUnJhx5OV
3eJX3If+p3qBzLgLZLMpOn61lBaJcdPT/dzH18tdE42IejsbaGjyZ+YlwRsXdIVk
vJF9UgSSf60U1PbUwrzRJizItTK3pXBBtbg3BfZaFyYgutqYJyddXTD7ngfKd1V5
LE4HAQqxt38JASWI1tTZ4PAjeIK1cHjr1DA5n8QQ1/2fxB3EcI+U+QZYFrghcCzx
PB9OT5fjIIEGJUZXkfNb5b+sQMmF4DCzn0z/LSRKMruIy7CRMqipK0KliIFpGBhX
OBfgnyGxvYzRntieeHu/cbjxjCNCpOf5jBU1zIyOah9T5/edboB75ylHylyFWOHo
2dJ5jKn2XgXbM4LOLLIM6DLZSIGhtg4M9LJFWNvTITXHi9+N5hIrlFjQ1xM5ZKXi
qh8bymVUVRfkKssyqWbqBd4donohEX7MKeLzjBviAP838gGHspd2/bZiO7MxdWbi
HD5krG9fSvPyNtFVGhSKLqNwTz0OAkE8obkb942jMH56bWGoj8TXtasSDiFtODwi
GNinWPUUna6hgkzLxSZdBnuQy5tWGCgyHkSbuaUP0NPJUGsR0UoQ2LeuvGkBB9Pf
gvjZf5tnr2gAUiqlvJdNw61B5+NJjuFGAxWPchRSRFITvnEMmEY4fwpsEh5gG96S
eyG95nFgjHN/6hnRM6IZYsZcMsf74SGhFKoEEYVk2mQ6XAC2wxrw0oqLH3JiC3q7
6KfFUvUY1A+n/xOnUlqcA1EPuMimd9aRn4rslzXCz3HIGaVEwm+P8s2nrSc7cKhd
oC+pNdAbv65ma1xVc/we5pksoj05W0mJfW1jzubu0mr7PulcJ3iLwr2sJ+ESOFi0
9jjPRi10ddbU1R4CcZ16LqvQu9t6UlFCAmL4FWhZxHWNeWqmnlJjCXaJp0yuJXpr
ZWc8CTbEiXWXOgbwwzrkVckv/JamfHglnmOPRsPUEJy91jyXw1yv5bsKE20sFu63
j7awv+q5q8PpgK8kUrzAqusgNG7sZNADN6OP/xCFU/Ra9ERpEHQcWzliXtbrodz2
F0RqGNr9khvkz3YGiqcwDUosYEK3C2DhIAj+PMcGRaMlDaVc07OXHh1u5ixmepRm
q81UF3d0JpcES6DQI6S6aygDY2rCvn59Ivo8gDveF86RsfcfK7PbB6xCo9mBxgrE
qubJBRpIjgZFlqxWpQP0bmPNUrr/jravPz6w+uufyumVaYN/WVDO7Af3ByyY3lrU
pBW9T3P7FcsdF3jNTJd9FjBU35ipuLfk9CZP4KnHZu/Wl7KZQPhxtNz2C/cQs+It
pTrIjSE8GEUa9gaRS5IaOxrQuDooBbgSoU5WRoYhmS53tUuC6KPyScmLH4ZpHwtY
AlYYKMcEtmW5/fLmFNSk/trwaI9e9PtZu4dKvDvrw6fJ+cXIDTNePl6k9NfF0hUY
GAQrspogQ/z/ba7NxHWN78oLruAvm+PSjcyy/CwKMovs8v/wj1WaBo0BHYeIPKKx
awbu//owXU6NKi4Xkf+eeKm06/k7wKuYDGp2zWyGOhkszkJTaIYpkgUOkUYmfY8X
6mD6vOl7EbOrPYNR7hQbFSkqagOXUQ1gBOo0VY6bluiFr8la/N9y06MTeXGVpoVE
si219XcABq2e0edVTSvKN/mAJbyRSEN4MBZctiGGULhBumwHJ4Z0/udgpSGDeMki
aIkmuswTzR8irw3YYHxEnsa/N78q9I4wv36YD7I+pKgp8xtgxOzb8w3GdVCo22kG
unr+35pyiQAwOjifIAI62xMtOQkB549tTXZtnjJvDpOw6IhF6oMu3ZnqNIcxf7s8
96HEXU+o2L02jm5jh8fdSojvrWLoaFKUjtaOv4AxhSOV7UYVbZuRrQSwbOr+oKxj
rxJG8bhUgVCuL6QAPWhF/dcrLiN+f71b0LjKOGgg5dKBT+NSqDvyeTJX1MrXaML0
5yEFXGuslufmSTdO8Bx/HPltmKOtQqTQBAn1uT1SQfpGVEyp5PfE0hPKDB5HPvdf
+TOhgVETylWDD6e2h+S01lskE/v+PGZUdUGMZcgv5Aqyi2FxzkEytQ35j5rztIO+
mnsOK9JjWiBRihh6AP135JVIXdYaQwlLmOjWiX6ERiI7tBDvQ8xxHcj14vs7xkMX
pE2qFBxANADsArR5iIGb9B8M597oqPg9OSDAS88Td001MtfJ6Q7aPfpOUPzM/y+1
RNonuXqm/F2MwRvthMf0/SihE1XeOQbpU79U1RvvcpXz51MI71R1clyg/6/nW9KX
/fUR/1nEBRESxr7dmr11itQBxmbYjxEyVNb84SSY2lOI0v1JT7ehDd5HhTk/mPGw
TlzmY5VG+E39egPhNILIzvrHMZrwUGfDueu7Vj2pTPIu90vfeHFBH3YyZ1utg4pa
kvUohfEkLeuAMljfRTqkbPR7sMPa93zSNL9DK7CPLl+F/n5c8ZIXFzl08RJfNm+x
rDXh1dmO6bUynRfrHO41gCenWD6fVSbsti3fCKiXw9ztjS+wlk1p/rJu+BJQ0fkR
wRyqeU63XOyw+p1nw+8bSivpnhFx5VrRbkmZ+Su0cqIJMY03e82bPUL9dIUbgsbn
BbvBujSWLJejlGQ7MqwDJUCCsGIoTGGVxtfclcoCRbCkN65DXUj9qhNSDtLGDiHu
lTAPzS49MAPUaLj3/lu/YxRsQzlQQTcnV6tsGcL37gEurG+oD99ZhJJCRmaOMYlY
I88olAeTov5lNkitFQ0OxWglJVT0hLkubUJM/CaDssKKZzUyrTk+exSvN+Vh/EqH
utf8cP/dCanpnaLa1rAR/5DS5DOQ0yxU4N0ur0WTKv7TObJzYX5XZGGvavQk8MHj
2c48kIpTCc0q3T5wngGd9nnlVAmLml3S5vtVR4F5iqs65lASN7M7z2qlu67EPi/3
fwkj+Vl/w50MLT91ivAdl1m/JXteXH2P4oSZ5bJaR15y45frEF+XFpNnG/mSuRMV
SDh50tdYNa8rjK/+6vLA5V2pKHWAeyO++6zOW2vtnb/iiawPSVxARlK/hnckeq2Q
kuPusaVV3+ef8O6AWw/ePql7xtcFK76NU2lDDhYqFwESmMoKTJYwT6Az12+++aW7
IzNrmB8htvSrqBwqenmj/GXTiM4Bpuahl/Atgs/BBkzGOAK+ZZ4n3I91EI/pneRe
Q6ROJoFEsrBqZjW+Goy9xzsLud7Q3Sya4jNckpiFz5JpTvsl975A+654wX0pjdYA
VAD///l+6eHSoXWfyz9VHMhfdlEWgN1MofE0Bhm1uBHFlYEkIWCB/LnMCDe5ZbW1
zbspl9r5nhloG5QRYryRVIITmMhkbs8dnD/jfqbjoCzHn1aDZPCiKOCE8DrkJSUL
aRoAQgZbyf/W3SPkI6eE5R5dsty+JzzZDxdhJF/M/0ojRHKCFjqN3EuOrrtHtnrT
VVwPPgR4PTkkJ8co+Vpkmt7ZsM3suBK+g4pqlkuoD/Vtci3My+SXRsaGoNUL3sNO
ZiITf9qYGuG1ilr/LIjaLK9UHReNOE2f7lXq1wz50pvCTCu18XiLoXanIGK+Oc5T
lN6DjLU7gdKIpPoASfETE/LQTwcdb54mnIM9H5NbsnEcoEyjvXHaOQ1+CgXrEWxs
fEePKZQDBV6u/iPQIU4StVAq2nothS5KgWINSn2AQP7+RLGeygriw7QHKbdRRGo2
HMBzOyQqae8TnUoknTz7I1l43S9Auo2lBw3VX4qJUWt4wCeHkrWdwHCSsh8w/xES
PoIBBU/O83VfxPIy2H10HVP9+7+IStxdj9e8YGiDOki9OCmmUJjiwYNopGMaIeMS
43RSMKp5U1V0xTHTf7/XPVNSPuozTX4+dA3dB0DAxBKDAUop4QFGpR5GDJ+IWy0X
7RJDC/YhixwKUfs9n9NGcM6Ire2LxDqFgNxa4IZ2tRDJgtjaJi3fDLCVJ/PyS6Mc
8/reMinAxnGmpO1wq3er+IVoSc5/GEf70axt11RO2QJjk1xwQGFSjbQszX61KyEp
UuL1ZfY8g2/DDSYPzYNdhoD4pLGrtDiFY/ARYQWm9QKUZahudu/4TgktzURZoJrb
0btgK/iMZl+pAsoWf2ty8+zoxiYSCvaYcOvRdmUiWA1i/18G+bZzUWRHbIklrAZc
qIyY0m8UABvjJLGey8lzrmLCuTXffhP2ZJQHqcsB6GSF886+owsXMzNnzjWN8pXR
yJIiO6sBMg6SOfTEoWYQhowpbj80DBYiiaVW9yTcixLdd4a3bZXHORm+4Fh2t7g2
5SAifOOD0xFjG9AIfuBQwgDOkwGAoCZWomc6BDgLgw6dXl9i1ovpWppba23OeQhf
dxf85nS9EssYHNYSxqyTqCZOEAY8E8lECjyGAhciLc5yPBxP2WxOusFFBjXP4VqZ
SvgvfLVNkyTZbZPejypXGbAgSsDZWYRQFveNjx0sq7EX1kwfvYXEZB5B6S0G8Ird
pHNd6O/r5c4aJRgRqRyBwhZ4qkI8VH3/I0MyPEKo0ZtyL0RTmWKGxfcB52AZu/od
6GoNelz2s2KWhacZlZY2T8lu00N0Ovo7eQzAE46v0HL81llWEqAzwy2iTTZxAlDp
vln6vFgcmStvAxEbAmJHDacOa7XSojOeRihhEcmsOgT3xpBUqgW8lPDKsrT9f3+I
qUJGvTt3TuBy4yVJ4MaquwmnLZrbhBgQn9efqJv16LeNXZuRtrL2wmTcoUFrd5md
3dgTys8IrLygoDVFbFAeVdnCuZyvWswTmOeRVlgdAYO17xqjJw4w8DaCWXT++vVh
nzLpWC6e1EFpJ5lilCjdtWdlOABN8xT3P/Qf5GOK+RWDkYEpEEsGbfuG4NTi9O5B
HfFQtlihHh5rgtLmZEHm3VS3lWwoK7xR5udSSjwQc7xpy2CJ3wejlq/xJwYVEYt/
iH72QsnDVuiUcGJDda446eWtVzOsc69d7omxO3l28anQtGnNcS/2l205wP9YLss3
yxuPiLx4nSAek9SU9Tu/9JQUFVm+i+t/m8ESZgFjXPuK3AlUDttB1i7RwFnMH3Y6
8O7gzRJTlPWIMRE4+F6yQb594eWyaw88nUS/M5h5tlS2rwU8IURO/Pt9KV65IXA7
xdWwlqx3DHQDJL0CTwOJgDmkVYpBRUWsjP7hpQVF+OG1ak7yn+AsImjkdhWe/ozX
D/Km/65fTQoACbyufy6XLEg7VfEkajgmgaAIIcNfMCMg8r/df5gItSjOxG6PIJdM
a2Gh73vzJBFbelmfhuflToq+P951Dtzk45PK92vXh4eBerHE99p3dgTEzmBxvQ2A
NSFODSMYcuj3D2kJuj5kVGsO7uI0c46Ls79sivWMYWPZ1rJJO+1V4rto1II9C1OH
sYOkiLqNTvPib5uO/5jhoQr/owBofZiginkhm2Qr6hTIQNTV40ug7wVen3OExhbt
p5ykKOxTVCdQKI8s1cKfLSyiBe7Io7Hb3k3EbzuACI6mclET3HLRODZ2KWypL7Tn
OxA8DdljkF2ZXOhoLVA3am0pnKUG8Mqp4GkclijXMSRcS1QfIeJ36NZVqD2aJ+Ci
VFS6aOqF59+pZJIPcKdla0OOabwIsx4zIrN1xDjvvr5Q07q+3ovOBKfTz7yUi2ap
MMS5fwyPXfVVvJTLRnuapumUe1+quQzQF2cW+FAj6pHOQ0JqOqo/l1rrgbuO/1ZB
i1Q7TANIYEKfW9zmemYu8YlvqZJ8TFPUsKQ5GxXBm2LnfCshZoZiX/H60EnuK+O/
30ohHdPf1bpvyhcsSqH98dnfSRxkszq+ySJLrYsivWgrVxqawRI0CTtsX3AcPTvk
6WXLHrKT2zlztwybHA99a+o9xkKP9PIHjkaB04dwu+QaGOGJK8oklKArLqdj1cRG
LRlTlZr5y3dl85haJ7DE2+DHm+5rTIE7WTJF3NNUyiMtcK8nLzvbpIALCQKU+D34
hmfO0TrTRfh/KL/oxeQ7DF8E8DMW4e+Fr4JC6MiHiXFwzB1w8VzJiHfggyb8gc+z
Gobp/QQlEuPujsQiANolFIi/eVcr8nHSFjFVoKOfouMMetfDPcKLXyNkVyuspZkn
oz62ZA9dVu15B9M+5g4T68xcjSX9Ut9QaRRU6HseCgbbLj1gcVReL7z9L9Lt0GxE
D+1sC4RQld8ULuln84pv50EWK1E98WFmEljSfD6DKlEkmt0qmu1JZpOqSvyziLiU
nDe6JdH0FOxlhnlSXiI6H480CeUxOzZ6/RQTsNY0wtxd8gNI4ngdVIDzyiGZt/71
qHP3WdH2SMjnxq7xaw5Zgijf22lKr3MFdnxEC94R7CzVISn20MN9NatAqHalFaKk
k+eEo/0g9hrlsGFTovWZKw1lgcpQXOXb67lINjO+trXO/Myx0noSNULosMIdxIi1
YDGtf9dbh9xsiYw1Ut6AlJjkUCkD/nc2TDK5qdlg1Gx83R9ocFpnn1gu4XI9eul6
6bdXqHxdj6d4qkiN2wayO2nON5hUNxkmR879EIf1AplaGFbC1graia5a7K+pQ+Ht
2d5RmIAq0DDiK3uHCm32+tdAOr79sRwbdN/mJ0NojPXW5aghdluWMf2+1TDNRoPf
7Lgp66nFwdNBVMZnyw2NjYSwKPn+dq2HR45x3fV+U3CpDVcGKa0FdQxI5Jlf1Tb/
8pWlI+MVY1ft/UwLTxoSEWYwi8PcgSxh3qMLSo8CDPjpgRpjPaE2621cYX2//J3A
qk2XW8adbsfTKE/cwdGY8mVF5i+/1LOFvOR31mvM/hKf8iY84cVY+ej+78rFftQ8
ZMSR76QOJi4vXBZXDQDzYOKVA46RSq67Z84+Z1MWFcI0eWJoLiFjYgNNPKDc+amf
PhCHvyg6Z/lmFDvCOMhoj8XW/ZrsQa2k9B8V/RjWJNplG/0xox6hIuGz8Mox4rER
sJ2tOa3r/1sx4MbiGR2U+/tzY9by9SCDsSjdCB7eYU4VdKRnZ+c9KcWG7VoG/Iv+
mlX4DyQiw1CFgJtMVF+BAKVwQcvgTpFHRP2av5CiRuMyX7uJ3YC2LeeUfRHLh1mu
opNzLpUfNH9oDdAvXL2Dr9RT9hBWtEFAGWR3o08MG4gZoncI0w3gcxVTqWg7qdHg
xIfbCqS7bxL9MrJJC86kD25/NDtank8DxKVNjn/Zc0UwbCnWKy+7hQAjWQbHGVag
1+4WqOLGz9dRcb6IYdB+SjA/p9zcdc2ZMMibivJNrKdNXsY7zZbxiu9wL5xXsUMz
ox27zPvDPsm1SCni7MQRv8lkufQb1z5pr2AZpxyGqq1lAxfk79Yl6krY6r4uZ8J2
7wrVu96Tm+snlxg5DBmL/631BCR0RNJ4oCSwd5BUf4LYKQV6GQIB8TcqcRDKseHT
+64Hwudeql2xq2+MsAQYUoPPduBuEuogeKlWt20553WJe74EtBoGhH5YNjeloD/x
9ICd4jGmR3e5eSElB4O1+Yl1BFqW4A6HxTdXLAnv4r+GAOmwwTMkudLBAlUjy/T0
aPUKIN3J3Id+z/chcJdkJdcm4uaWfWWvbvd55agQoK+ZXybuis4oE//xs7D6LRYl
vf7mHgtoU4eLRjAYOYGDOz8b++Gyyho1zr/Ruly1dyQFaTEA69BHwmfBtLk+5FF2
SuAem2oBqXtbRMI0hGbmcI+fgctcvxfi2TzdB03zni/6yNTXXsTysrR71gyykdOD
L+mtlCfvRRTKNCDp26PSpGNO5FnTfChJf2l1XOaqMhucLfa7RKsCYbWRGFnxcci3
gCB5kezTLPTsBmPn7iN9r8J1HJ4jrP6+NPuNQ+s0EPoElPjCByMFFgekempS4Mxs
7SiJH2k0gOmKlj9Yo5qxlQlnJZ/01nczWqBiV3eaoMCcZqbV82uHhgCftB9aujpx
q8jjT96gV9cyF8bauO/BkxBmn7NK8tbMNqT8DijmFAWD8K2UcG1YxrWi51AxpLHf
W4KUPGiCAtjHn/IuWTZJdW6Gulymb1cqT+U/Iq26Gxzdss7NupqPKajJeK/dhd2v
yNLmAfGVo+IeAakH7KOsDxwm6RlO8Mcac2bFu1wHHWcQoETaccR5wyNEqRxFFoMh
QaNfxtVqlRQnyj3gXB3Uiia5gdnQyg8i0A9AUe29SDmd8sWNOO4AKQFlGm5VZtej
YW36L3Wym1dkvxy1TP3/l4p7JA914b8CDoxS00Er/0BoXWjhMKGAI6DzGfOWbWq2
XCRXL9bzD+G9G1R5SbHfFd2ij7FLNH5yzrI+2rbytP2TEV6UGA2SGYv2hEhU53pU
I7g/CouOKeV3K1letwRGeVZEjbibKJHgT6WKDt1zxNEjVbl2M/QSaMDNNlw3QgwZ
vz5jwFZKor4U85pwh8NPBp87TqNQj41OA37fgTfaHciGBnv9FA5FvFXggD9HaDqK
8+koGpSLy4GitNDO/Ytg+3zdeURnzczwQFlb0pwBPqtEG9yrEYw6tI8hNT56HwS2
tdwlRTM6nDsIQzsWf0Yo4J881ns/CVouRNnj8PJsrDcAzr/xyYoro12IIckmlWzC
GEXpnjpq4oCD2U/pqenU6lk5EDOvVHHEa+tUXWckbPED+Iy6eC/qFj+am91ZVfM7
+mR5iWvG/4Hn6TBRkWb4nt15FwS8K3O0FNuG2p8wmifpIQ6jyfbFREFAcgWhuzQb
gvJ98EEIWNka44jaeKXoJDAfSTM9EG0YXjx30Fn6fV4aXHypUr130ESENQ+Y95xe
KIPoobEmJBRC670t4dC/0p1Vau9RrKGd94jrLJUhsHaZ0jg4TO2oF4/nxnq075fB
GO2WCGSZHmk8zvYWNnQ7JituQjtf/jqJPEsfzF8ysQFknx5vuvlMMQNNivBXB7DR
IN8FM/GJlfB1LgK5G/8oJf66H6zMtxxRHzp6v+TJe8Hzkw6XxjRXweowQHQWtrDs
rM+kVtra8CDbLMR/xeetjl4tBGMKHzx9TK/wPRa/sMHJuiN0lXQEpPrBY9gVNNbU
BkqCkHVwm5Qe5Ma8/p0Y6cG5M+P4hR+m4/UmyhAthx/ZkqRRCWOLq0PdOYWCYCzk
eHQLpUiay/iqvUIDD0dh1Fv0Wme9ztZLV0Y8SEx+0SdCKOId+W1HAOPpghekbGi0
mZLqcx/5bHMVv9QfjWdB1SruEZvZKnZv1RMGoAN4yYtYWQzfI2HSYlmd0t10lvwM
54Nmsnkmy9rIRqbCjTZ64x+xtnd2l0dFz4giztO6JHo8EaxhzEzzI3YvpLz0URdQ
zpiKjs4r26FIUoKxbFv4p60OLt+525rvVwusps8VoakLzgQAclL2JJgR3LuOR2zE
T/ac37/8wK+ITfHON2kRyARBmEEkPcqEzJIuo7Q2ebDKs8G0WFoaaSZhjkz2M9gE
N+rF0SMhKmD+G7AalaUXIhsKsNaG0gbjho/rZhuVif5CzGErBFeuGiob7UB04w8K
XtwqJSntiI1HqWEiMkmAmKACShI5YtE83AZ6HyT66FmjPy+emWrGC8YdPLjnuqJ3
8ENBEKWBGuCJ8h4amYk98buwafgjMvDryziwg2j0v+KDngafUtcZvQDWurzbpA8i
zELUYrZFRpgJgbWcwUPfk47VBmLlHOLpcpuwOwFhXPGkzW/oNu7p+/7qPoYDIQcQ
GRTxWm7cqldgJO2ZBGzOiJjuF+3KUOvW5VXykZZjlMYiMbGdi4+N6mTYlG+iU8jL
xWNQieTxKXjY6nRVySs95YVYG0SzmHLq1xiUjHJ6/siz7zZOi3v/qAYjG3HG8LJp
GRJoMaLglYbtEtQCuqY97MeMbBNCInwELJaB9Xt9DUZZ1B6uh02YEgMnh4tkskGi
5PDEU3dbHedqa0uJUosMHn00T+ChWuI6SzOEt4E6bx9ic09dG5rSJpCN/7Kc41Z6
BN+zCh1aBbWIMPBUrtcPjn3ZU08/tJyPIXScmM4fJrWZTOaizO3C6mDNMHzTpv9O
jm1QdwOZMqNP/RtoSE5mUw/ZS8F4tsZyF5YMJ5K7HKTAeejvn+b6E5wh/UdJjrsz
lpXu1twJc4c6YSAkcXlStZwP2Hf4lFUiPcaWJPy3p+LfKLffoNibpL7tJd0TJoJD
AnW62sCfRhb02NzUzdvv6Eq/uAFErO2POSnH5BLRYIBSRTGcxpsY35IgzFI/5az5
Zrxbk97pVLr11QJiXuhBSMG2cjPQiF6AGhQkzMEId61isrPmdGsi1U9oIy+gSf6v
US9qVaLmcYNrs0xVEhorxuqnxD3r4xQHMutdMomyQ1AjNaO+cPH0McN3Y2kRtzXR
grz7ROQ+1cejR3pK5o0K2FRnKd5Adda5uHQziM9D5uiRtMflUJNDj59tCrdEWlkt
F30hiSNbb/uB4FIZ3HcMUz5JibApigrrRQIccanfFFvx9yUHwrgy9MooLcfnsHPm
b7xfbgHO845YJgKqCWmpLzwrDPeix/58Z4J6FyGcEm8G5+9J0+WKjERPQZ7/DCf0
JdRYBolpvO+R5JrSMTHVDzl7l13rdSNhTdB3rTRnUzai5f4WVK3j9myuRWfcmkuU
vee0sYQE45JPXmdunpacoeRKD6Hv9/KEVJinHNXJuvBORQOQI7vEH4FQrUlwa75+
UluVpxm3eiWBQIgDinu7txOY/YozDPyGhWxzyt7guHAE/B28vpQaVqJXPb3YEBYn
z4Z0DkHIy6cHO/Qwgij6UUk329P/k8YARduS1QNY+dJxzAze5KTTUCufK8wC118a
Sgao/PnhyqUltPMpiJhXN/5nv6xdjfUUh9j8TpAXHDhYEQRTh1n2jcJGF/ciqpkQ
NdWVAUmiCc7czSsx87VUsxIC+w/k8w48e+ctVMqrOhR0zgeaqrHVyAqYcTLOGyzu
QpIL6fMplcnVIIEtohCsPDiybDaOSqZrqUrYjppzqFsm8SzuXnrEUQ3B0OdCM8MB
P+w6gySwB0HpLvJ9yUpCF6XAad0XzLhhlZUWcxlOwKEhBmZmivhsM9ABe3es/pm1
zzcEShHWqfwcWIH+75DDwAUZAj4/El2XAS4jP2Mcr+q8hATyb2Va0uXI0CikKKaW
xfM1G3KNMai1OM9vY4+B6MvxYkQawqQi8ZV2wiihenAKOPdiIrMSE+h34Z4O32mW
zrzeuJavqCWNSUYJp6HeNQC5OogmENw9KBuVq/Qyp+jv4atU5iGj0ODwmHXz9Z1R
2gNtlXEG5/FRyaUQO9uJso+bD1heW5/cbtFlyQ3Gnqu7Nc5i3uqVFSevdtNVnm9b
YwL2A8cvBzDzUBo/rTFeVAITISgGSbm8Ze/1xKwqfdEyUApfOEB4VHli6104fTfc
vyDtppKvF1I3Ma4Oib47cOGOZZbPr1I0o6oJPy3gYLdLjWD2yypDcmcp7+SVY1CZ
+g8FpWj+4UhveN+aWIpnBry8fnIyRHWjv8z3FXduJUDJ/gm3cktMsfzGD+c03oIi
mu5fGM91CbgB0E9qpyzIbrsHJ4UeNoo7HbTUgnhDU32yPkQSkz9XSjX/iIOgvUbA
86UcKrHg3370e6QSyZ0elwV9lj2KFLyxGpaXgqfLCK44bKJb0FY5TlvCTBfHitr0
AXVFDVVpO05IdJl4hUtLMzCF4Tg2Q9B+xkhsnX5BAGOuZSKby584vPcB6ThPnTQ/
5dSf3LFHFHqsy4lG5jUYeR4IEXGbWz8HJN9vYPtL5XdOQlvzVchHcJpVQDiod/J0
4SDZwqaUncfKZkbef+aIt1P6sP2o8TR3cCoY9GRjV25w1eOKFMw9s3L9QXaaazBC
++Zx/VpcOG39DGVIJND+yuPQgKtyGt5Ayq3jBeVaDY2pgDWacmDhNyaXTEqQpHak
wUAHuaKvUvd9ZgPvwQqASkTFqLrqarL7uaR5ooiWxBh1ud8JJ5tEn8qUi0HoteQB
hAAGMvywGr45tHdza3gqit50cKjHulQOAfsntFc1EacTQrkmxVU7ETk1PJVM8Ggq
tweLi6nNxRwNudJUoflJ0aHhfpmZj0+Tlm+ugBmsJku91ofXleYvWxewfpnA5JTi
tRgQLKol7gkDg7U65FMBrY4LpcUJVIXHUVq1AfpTuwRxyzpOSAGelW5JLDgYpd7T
fBRvngW2wSrNYHyhtAY2VemHH1ZjvWjWB2QZdAluT2/T/p3QRJbj8b27IDejuHGr
4Df7jChu2h/eaSl9V4ZAjCuFWJ8eL8Bv38xE2qbNp8fgMyWPgNMV7xGszqy1tIVR
+m5KCvNzrasRV8YD1zaryGbrY6aDnghlTlF/nkxJIPjBsHHhXZvLxBe0xhQLV4gu
K9yD/C44X2LBKUHB0pbuXZKWIJPXbpHHrhJedxAfxT6JqHrgqGSjzp1yvaufNVIa
ovrlb+zDRYJF53td+Olg+JRTEJqGhFMybxcplwPvyQYVaW9xVUkGDMiv779JtC3j
F0SErBDh2ss/lNp/UrXae6hAsMHP22kwfCmblWbkBUHIfakhw9zGi1HXqrXTCfdx
ecAvHcE4WX/xkzhNs70PlYmgFyrjXhUpyAaZ0On6XuoyOD5CEXx8uuVNcjTHPKBg
Ti7JejCJESbJNlZMl/EsWhNOXYWV1Sq965INYAGUtUawUIAe3bzzabSMw8WGssrQ
g4cewOIcv0JFbm0Jl8deRfxl/1buG+pZNlXwcgHYdvGpSzNhk+1TbI9zuaNrN+jV
zpBXN8eXY1CcUrUlCF8VcC5c+tcuOpVWs+0HYZCVm1hxZXBMFDdDM//2nO8cVlZT
26IK7TgOB6MBb2W+Y30W9TyRDlJ8AT4tjTs/6JSgzbl3yCupa1mEC24V7KXR19UQ
ryvumNcq+4nZue+5tyM+/XCfIlQ5g90YzZS01P2TQtQlt6395TpgZGV203c+B4WU
SYx/VehiD+6vYcIr3yWYINFLATnmlwqJ4iphE/eLnJPX4prr86I3iQ3h7QBA2M5O
JL+DbqdlUPbe9o8GFl/0YQudh5HLYMFRUS5x1lU0iHgi3ZXU7Aou2zhix3L8Mua0
x+kf4o18y9yESbYrlOUo0XA87K0r3T0zUmSBx2Saf8in19BmNP07pYwvcR41uo1f
CsqSfyCjkMl73ezUYyqtxcFgo4dkKrN5qmRYZILyeVthZ5DvVmuyacaHZzbVz3Q8
S/n4BUNN73EQVkSh16KLVAdj+wp+pIzHp+wK+wVaRMy/5VAyw4LmzF0VlUC5Mqn5
c3z+GPm6Hn/AVb0JU3DYwALL+KbOsLb/9t91WQlcPC/RAEJvohvdrzjwtJXoxFOf
5/rj6n0dHWAAoqT2AXCmqlqclN3GhXjZGegfhTrT4LhBfen5L83gGN9FbJIyOzZQ
HyotSmyW4cY2POmrEuYYxButXUIr894tIAv8Unsb2/8rHC/NxfEaB+I9Rc9ljM2B
NAx0HKXUeG6IzURJZuHo72X5m2HLGODUvuSfbpnnpsKFz8vUUSUfPTPD1ZLj6bXN
rOzryYBjGopsLoRX9OpvzQXzpDeZn7VNFAjiH7e9+hpogl51d0KysSuc7V25r1Ep
nKAkgML+/q0NZCob1f4EDnA2/g8YYpBEqQFEH8W+t+IzAU88V9ydtuxmtEwevpT5
UKiCjvMdt9jiy0N+Dx6FuSecVBMzXrhj3FCU6WepxyCaRJsJtttLJCQIJUxRS00h
r+YQPOaTyBCW9oVrOqGSO5RWmRj2dkp72X227KZQA0Zp8xYEIQtf1TY8seWelVhJ
ewp/FkZR4Pw2fNKwhJumlrkBroF+EmxanT9igyQgs0WnaFmchvpmzSsljYFEhDFh
dT75pI5pTbtgGCqCMoswYQMSG/Q0znSgqZyInapuEq2Lvxkf5wBK7Tan30PCuf5o
J4c0LauZFiae83XCUV3mF/M8ToONoaT7Qt55/Zf3PZCDxP532sF/1jf8kSSaK50X
oaudSh0oOVU51D8rpf7rAaPja+tS31sy9EqPLTdfQvtboCJ7lc6KK9E7cyw6NKUI
pHJMLYZm3ue2wyJgWPRASAl/PHLtMrolt8yI8HXABkWLHqefiQ5GaOBs5jV55LG+
QMeuitNLHKmGQ+wZnA0ywP/fS10zj7uqKdL980zaPBkbTPPUVjr4XLeTlVjk+9sk
193azfuLfpxy7aO/Lyr0QD4QPtJeYZkZWd1ZLhIFXi0O8y0otKEgr15v9GrZ0yp+
AJ9dYPphZL0Z7LR8Enk5ltKobom1an4cmr7+nQHKv4s7yfa2spCojRIg5wAmCdiS
at0sdSHO7WE1itAvZJnuRH8dtiMgLIahf/pzoHADfsp8CpqZNgBZdxfaHBWWd0Vc
INPvLNNJHNTprVauKQ1hZfCvj6EyZmJ9gHrS0D6hMu4Gyp0DtluIFjcOtGxpv4Ng
WYeSG17MsZRXEpWYJyqCHCLSwmmSZT3/3DirJvjGl15ibp8Yu7cvpAtFHwbDPU4l
q3VpAfchIG4rEtcuTcQZQAn+ZNuENf3V3zpoF5OZMkiM8Z+QxqzPxGFUCv/r35Ty
LmxvwTsQpDtoeJuVuaoc6Hjw9uTUdWLtwGcF1BS3u8i9UeWotdNSU98Spa6UrDdy
J3BAt5bm/piyhKY/0ZbeCicI3lC0LGNYBxFAF2FJkEoYhC+QrOgl+30gkWLs1qi0
/daH1JWficbNFp9qIOXj9qoAPiaTh0hkQp67F7PEw23XyqN2vuhmok147nOB2i1m
B3NKPaxte/VHzXq4Z0LWAwj0bld3UGfYZzbyONfbo/GcLP0R7jTP+Avfrkjw0ykF
QRTyqjc1giB2iw12m8isgUcpEFEnGFmQfYY7CedXy/ieBxSYajuKYDFM/GBKIYlX
OkULWkaqU4nXf2voJjxXbhBwX8w7Aj6s59+9YUCdZGn6nnvAT9fQ9tH6LJLUICVG
EpP2K36qnhzm57JZ8FBMk4f14Mi+7kZYWyXIFTgoY2nNqux2dBsccEZ7GfiF7uh+
JzWqyP6OmIeKu0baXxbTdIEktpS0nit0vN81EoUdCwLX232VmpXdWhwNrc1QuxLl
XSN6z8M2mgEhtP31NkoVquOPXVWaCHw56L5C7p5TLsedAnqxBuWgDyZRJz4lz8FB
/9hJIvmIYDbRqpKhh3K4ia11sAcJfJDvi6dQElD2yYb40RnuoqAzKl5ouirW+rkC
jdAaPmmvE5LV3xw9zoGKQfh/QLOvLpYsbltToEewrSLN00rXyTKk62Kq8NlQtYuq
6QhsuXE4+mm6/2JwD/F57s227eCNHnbDdlN4tBTpEMOrGS3KOVpAGtqMo7Y2rbCm
wyiA8pBnXw+9vOzFAvC2iJ3Q1CuKnnJdSw9YAahSj4NgBPBOipRmNr7xolGMlxO3
YYtfqrr7zl4OhPmzLP5jtcOOwLKGRV9uCu2D8K0bSCLzGPjCZUvGh6XW3FktO8sF
nPc/Vorg/H2DEOxniaJthNtf5VtcRJa/NzZDp/jSUlZT3th75Er6gf1fZUtsSLR2
LOQ7TT1/U7Wg4NTTLD32eXtiEaLxRO4Ga1raLH8t1jjPXG73Lby4yO17T89Pxz3p
xdsIbosqT7HM9+tcT0tksPjKLgcIaR4hgNFwb0k3wm9ISMuQIMysu4rfECp5ZAd+
V89JZxhKvEaUdHLHqXgMFLcHI9lqK38cz6Ti7cgjVG9ew71M1652U1cDynrYMj6L
HnHTYCRv8mum0xl6h4JHuALbJ+TST/hJ511RfVIhXF9UkxVt8RRKvgX6NJjM9elv
NrjuPvVbuU6fPXH93slKxsI9kwhzs2gmTGbVmMLVYaJ4qq+VBpXoqoZ7aWfxBQhD
IY8oxVqXdM6P0CUpI6EgVfnlBMNutmqJkw9WS81gm8b8X04A6O6+SXIjqkNqThfU
DJO+jN29byqLBB8luwLoAR5fBwINDhDrQoIADcFnU9nUPkYWLt+Ujncn0h1EwmHe
V+CMQfZr55tscwYSTi4qAUWbvlpDMjT8OO8kZ7frmCuoIIqEmpDFsG1Kg9QWQdzn
W1pa84bvrdSTSekPPPiHjPqsjtHJLq/bmXTUCrL97BP28L14lraUXPXsLa1me0Ra
XrhlrKiBce8XQFaV8UAOpcwGbQApcrqsEZMN10uem4Ep97QfMGmDxudpLV4LxLpf
JVd1zIO0FuZcR0d/UQQ7I4T+R0ttLP8BgeNP1Ftthmu8NDrtDLzOk228DsoL8mss
Czu6vU2l9hnTvS9VG9GraDVwhR/hOceDrTM2MBGtTsg6njt535QtEduH4tBEoRyI
YZKuG/pjX7sDGrwVXKk/5xTS9m8mOm8COco9IXnT9px1WRIFzk9JI2qUK+ixvJg6
yPWEwhF7deCxkwgu06sz8Y9KpGab0n73pKuSAN2ltgGUWh4uTeEdXdCCQoyZnYGq
8xzFBJlDB+ipPJLv3BKwKtv8qYaAOH5WS1sCYNWp9JlJp2GxOkHBeLODB8nQixBa
xcHq4ePoC07anfqrjFog4NZQyilyRbGq2LdHvh/vsdtnf/rMHG2nSJ0EjX5QaxFw
EHfKxz9oWrQOcQvt62WnE7p48ww6VvWCz3rcc8xZVg34SnFLyJGXDXUEJQMRDAeP
nF6/RxgCwlt909Jp64Gy9BB4cShQVsxRfLR4FKP/rbKa3vU+7WVBz5OxQr85mxND
EGn3/L7KKWY/d2F4xWmnHEKi6tuJKBQQlcR34g+UAT3sNoPC2c/6Z0gtd3pMKSFO
xxHhuuRTDZeUX+F2uR9oL9aLz717CUWEXc1lSRjPjTmp9KIxBPMy6nMhsxhtcDc+
vXwQCvtK+plIdSl39ME29D7RdHd/BnNWcFaI9RF5of1SXmYAl1VGGb2gKe7p1Js+
LNYFDP7ZwY/mHCZna4o8jBn6g65Suz0/en5VXYa2rCT2UOffSlTXf8JZb9mZOuAW
/W7Nea8zH9vk4fIyCGllyn+pPOspwawJ3CQWAf/7CZ7mZuVEdM4fplGb/boXtw4s
3aBgQGKxaGl2yZTn8Pkgu/SIHNWB3f7bdhDEr7LQTwn7aM16U2uCVOyHReOmxH8i
gKJFP84kLyCNOsuMUnia/IvbGXUHwEIEd5CugO9B1cYKk8MEQEavm4UtILVe9Imn
cu2nui0IO7G5mKGQu2ttT++VESGjT3mkDBJk6NCnYIzNuqDNAmPlM24oVkpQEbfy
NZH0bUQDySveYnmt+UIJn6J9auwWNfYUBWPmuwwkuWNJSLhOuUx/iXjibcbh4v8Z
nQbps7Ev8qjE74QG7YofdM5N7o3hlzG34JVIvbu1B9X5Okg6EPDcRYS1pJd9UCWO
sR72QQd0fRSe0lrNG27/pn3HKhoPrYBFWE31G4lcTKcPr4ine78Ze/ogn25nJxYL
SKGAWuy0QMT2a41N2mQXaIMFCo3jyg6ajpvDc0F360uglG1mXP6KXlaqXnAF96oG
AyE/7p2Tard8UHAph3CSm0ot+MI3Tt4nJx73sGUkUwaNvaXMOMWZQzwlOTyCkpDE
VODY/zjFOp4YR9Xbfj+mMFAXpELjD0Zu4fK9aKzEt8KacxX4QfLzicrTjSiaUv3G
BtZUxXgEqqSx8fOkTRr4G4qkr1XgYeA8OAHvmMNHbOSvRj9a3rH5VLq2lDnIgQKR
O2GkznMpkqViTibfZuhQMYQUCoxBBGhBOqGrv+K6kW3mnT8KYJMPJ2h2uXoXuXrO
wdRtn8a52iIJ7qspptG4F3XuLaXA9XO8F/PYwfNWxOiHk2rJJrK/87G+5EtP4CIM
pCbxyy37IIlU01m8XP30jwLzQ+Bnt8C5iFK4hLqV5HiiDwjMLCmy4ANWJmeWlAy8
ixWvZqpBehmmP1HseESlQp3zKp6a5inYW+DYhKBb6Q+Cgt/KbYmsdyn8+vc/9cuX
AGLBYvI5JCGLNe4Bd6XEvKXSG3ebkasi93V8tRPONh0jNSbzoDaa7fPOc9ufX1oP
TNu+UNnV4EEChNsY2TAlZceExXICcu8eiZxW7msWdYnZI/7SO0q7daBr6elPs4ar
uPZ6jGdd6saF3lwAsLUyfwbhBUb1lyd1UuFyqWMAGjrXT0wxNjaoolsboXAYubNZ
t5wF/1GKn/23KG+EpdPP47Tpb2yoDHGpLVYGhplrP334TF6qb1BiBqE6nZPZubX+
7XeVAAF25NmQjwGBam/PprwuBI5l/ynHWDKWGqODyE4SO84Jk5EJTJhiK7O0aM4j
Ku9WbnWGyJ/77VACEJNsO1grA4jbyKM47+pe+DbpuZvIfIQf0W3QY188cgIIiwQ2
eFe/J03ABKiic0W+9rflTH1ZgXgc5TL99ZtcclMXSwF53DUhfmIq/ok5IA4bPlX9
QJH+BieE5OYVK8QRO+0UWHQLE/RxhK59DC+AHXVAgNl/FaXxyyUbBb5QB155Mp7H
2YVWENgc5zbvEfkjhYp3fvNh2a8HQd3WQNltM41IL5Sfa+ZUDL0m/hrFWpk2pUrq
Hp9K+Z+qfD88Qg/57d2bRy0hbKs6T+w7eLctmzO37cP2Lh2dfSubdtmmK9BqPPw/
8PTjPY1X7WoPnmwix+/NRUJFVdBDVnUTpZpzqXNbRN5i2Rbv4PA/B9NpUSNrud89
HremBegq49lFXUh/QJVa01PkPcC9NLQM5f0ZKhPcKdO+v2VkeY06NUU8GPDT4cJ0
VudlioeKKNxI6byRQ6qdVmU2Q8aFLLz38yEHN4mgemqQPVB2ZVQOvYEKkVPjFydp
UYagJk3TBX6zuXUc+F8Ml+rU4Bsc3nBfENOTn67BjlVkApIWoPyFKCVMd+9ip5ni
zSke3h/zhnOgU22xLrhoX5eeGfZlqxZRPWbQKGSH9omX2lo21ujCurkMX+2QJfp0
Irpb6SJ9Jl8+aZvP+Xcl53yDfDngUO6bcySzmgRdAEqk7Bs754ysTPGO6ZOYWfEh
GrMwPbU+TVZ+wEVgmU38w8+k96pj/yHAxc1DB3AndjI5RIlXYi+sIfX78nVGf+qD
AbRSrf8fE3TP/1Ej/ev7/g76vbc34EOmpB6S40D5cEZrnxKBjrGt9SAu3M2Dk5x/
MsrruHHjVbKwn7yAYOVkYR73esh944C/bAXDbYUeiI9xnruFUjKgdpbbA271zkg3
+KZiTTOqHPomCsiUlFLlphR/N5c7mNlEVGA7f3WVSPqKfBYvps/ub8XyTBLbz/pd
cSTA5B7I+Zsf/Ln+Jo9ON7Pvm8/aVWkh0aG6tF8bUFRj95he32MnhxBCJ9AOItap
O/NWSw6AGdnZct5w1pGRkGsqMpGjBnK1gKNMyh170LmETPtOuZJ3pRxboRR7IbT1
86JeJmWwrMzz5KIt3zXqkHdpSRn9vDYCJ3rTKHFaoH9ahW+Smn48nPF2BRsVxxXg
eVV4bUl+pX1/9JGdjd9EAfsmk+ZBnuRKxrhJTFVVFdCltdyQoj5spp66e6sYCn9x
RSZcXU2RIUDrVUyCUCm2FT9+jyAOwmhRJzyqO97CAl/br//Osg0EQu2tc6fdnqg7
5r5uTjm1jX+MmK5Wn9yc9bZ6yqG4yuARHDdmta7K2jzmWdMCaRhd+mmlHOzsx5+6
Jkqca4VzPH4A1RXy1GEcxQes8xCQdFqfSneYEk13qwrxIIpoT3ZjysixZ8XHMSuL
hMPOfFU8cjebOfBcObnmoMQePus4K+7N+qR+0rhpev/mnghg1vMFKvRyqnZS2SPA
xODaQVzPSoBJ5thf7dZtH1VeAeJ2bE78gJMoUPm2KxGupnJkuo+kkXhxb/TkxJQZ
IdbA1qVKtc+Cp+8dOdGNl7sFBNXCTDP3vbJkvTXlnJkWav1UQsEd/E3i265/3z8Y
j0lxqkPWovV9HKR/8hMPgDx9jtvTWqRLFA2A4DYZi3avhM1BdhtFX6Bon82YWgMH
bfNwLFIDtY/5w3iSHM01+X0+lwH7N1J5K+TaRAQB239eC59XoTrfwmSEQlCMiMAt
LN0+tWcAEOzyuhUfmqpXa1hmcM6TYiduvnnuX1W3WVHamtNhbedvFmKZXVaiC54g
614VAj1uAZYUbbVpRqSy4nZffGPb64z3wOak9Jez1Cbye/0E31tdRPcEomvJYh/Q
Wb1ROWG6KKVs9frWejJZ1hnRI3GnpVmurlFp6ukeuCSt8+vYa1V9WkzSPMTZXLxT
QYh5eUbiLf20MmpopZUFLn/DW+mTkgCy1SEdTpnejysT+t/Kee1341INu3MUykLh
k5PARsGG6A/v3DByve71YbAxHIn0pMddNQdEiiJImu8S1TXm67XLEr65/3TtaQPX
jKsUNkg859ocKt2ZrdKmwfOqqOOjGJnQdDwIQ1HPhXYTPqNLd4V0nEj9DsuV4j5q
GTkOMLJpxRv7G4ivNkVFo3NeWG0oLJwHXkkRApEPZPoVbMSbM7JRpIZrGILFUOaH
iFeHZFF878yJ5wOGrkaslkX0tT72BdZnSS+3owtd51fGsbzSClHCQot516JP5wIn
KyxdvRk3WvIacQYtLgFG8k5mI+ZQnDevDgP13OW6lR1Pe62d/q2LSovwdryfTmeA
XEsE7Tg1p80A34oJWOH8GW36HNukxB0gfTvLIIRE9fAAtX4RdIRthekeKfogaOvJ
5ktqyHHjRGS+A41zLWAKoInwcp3vVvp6UsLGR4Nb6Gi4/p4Jj/Dhh4aQFIxlURK3
A9OFPrFvXZqT12XUkgs/k3SlrNGkIhLm1IIQ1oX3d0Ss+7+eavJQLI96W3USMG0m
FnKtog5QlBWKwmFGQ4ApfJMczB9whVV0czGO/M/qxds4wIPlPLpr6jIYIRTQM7qe
qyd/9l4r/SkhPUB9cgWAOrybeAvdQD2fn9TQi+chLXuEVexpC/GBz4dGlPv20MSs
W4XC+lMeBUPtmySadoIzjzKmvCdSZMOaj42YsAdGG73ynHmfW4u4u1ypp0grUPfX
68nV3DzhMpedPHxaE/6AEHCQk93zFAJHoXOFc2j8/XcR1+ip3aMSibmjiRtlSkl6
aqqK6EWFW+IzL8PVhELOV2g5fJk+XlG6dOnVLecjlqRacyywWE2oGEeNBV+AYl9v
W6UNKi7HlVHz81shCNlep0Ycn84avQepZenY7IfLwiQ8uIB3wpuS5F+w4D6xRtZI
caG/2+2i4ImOqbYf4oP2XDpjdmCAL6MQ0tx/zlizrWXGRovBKsVzoF4JnRd9P4iu
d2Ok5elmP8u2kFXOxlPZ9SfYlBDWLvJu4ydTFjD9/fbdGdU0c7F3P57Fwyga2xAx
PXytAPReaC3XuNKNb4KQ7Hz0CF1oUHYLJf3mPoai+ZbgPZ5fjjeLAtNjpZM0NrIl
HlPirh3BguNP+JNZOx1eWhi/ZHWfwUbeRUxBXd4EMku8lbSBXXihtZoT2P9xyGt4
S98vRDNVZtHjeuS7vKLKGRACxMnFiGvJVJdrcitU0r+tiNlhSiTIYTS5a/cQEs2o
8qUhQ8pZ5a+okOdqPHHaay/f6FL4ix9qHqzRIgIcXM2YJuYaAANzl23Jl7ZCGqia
Nvv7U6H1CeVrRCS8/kmRrNjJtuF9Wx1hQhhJ1ukGdvLV7BbudTwl7fV5f0IWeM7/
eihrdrNffSU8OHOOWgE3KLFUWIn0zpnQX18r4F4dW4AR3dwGC92QHyHQHnedD3Vo
3FTGTYKRXrcthN36e1iKERv1hP2fECDM9nnDW32LNpnVWwvnd8r+oudsvmAKVSj/
9qPIvMVUvCNv5witNLl2Q4uwrvxSROkqlh7pyJnTzMi8h5PDFwaGQb4BBnlZBp6e
NmO4U91fmXf5ahgD8c95GFv8iodfXubGh+QegOIaopUaXciwQMlXkW1+G0JB676o
ZgCvzLCNR1gw7GN+drrj48iBsvqegYUoMxYc5EoqWCTE3wOoo4aE01huzO9NKQhn
GR8vLi/k9VwqBewipDmjfqLgcgh/l4SS2k0f+zxSCHXWEn1Kzf3HRJnDpnkEoNrh
96RAl9M5WlBKQJXOi6n7h/fBPkJf+BcDDHdsCfGEn9Fi9dpwMismsCQtRkumqrOe
WFvY+M/VBSBsWt78XbnSacJHv2qtuv2YOP7TLPzNpYF92wSeurxxn1kIOVDm/Ksk
7IuEXTKCbAlU1r64ZWw6VA+Tpt+QfawaSW2Ut77GLlS1ny7eSrUPZAuIy0RhH8vl
R8sAw9nTDT2HIrdJTUGvDPzr8+YQayXYTZAKasokd7R+cYUPTJZDjiRw+Glf1faW
zry4KZXsXhW5zHREw0aKZftwJWtEhIgAfj7m4JWVlYAyZk2P5XaW3CWNL35wFG1w
sbY9/Nx5rnqKf8MHiR0jSNUmWa9VJNsIZZuNBYTLsgh2JJMgUOEIqpjD7YzgQjL3
uosEdxSDLFvhg0DW7tK/pEdemBLpQwL9OHQ4/0Y6FKc1DM0xO75yq8BHvMp46Ml8
OYkeFJwB6HfpUW7mG4pJQ3yoO9kE2jvO184RWmw3XTxJIjm7IS/VNLuGTkZ+vuKS
NEHvAL+esq4tvzlFd7g/8i5rCFojtEOdRTrMsg/lWyCTgStoI/WPl8juc/ghFczz
cGBpZ3sqgR14AgczantshAvYDp2y7R5FA0gXS4+yhk3wQc6KboJIof4xsh1Rh+kY
MrQqOJe4eGlUrq7wil88tHcGo9r0KNI5MIYcFeSezguOfQFdLiQXpiGz5g8ZBfoj
eWm/CCNxy9J1TRyxJEqQHgzpaWltso2CkVf86YniOXzkzx6S5DvtaZbghrwYthUf
RyXALKd9XkoOSPf3J1RUSQKcLpfnDuHql3YxTSu3I++a3MmRnyGZLM4O9klO4Z0e
H77a4D9OyIyMsRm3rcBHwdNnZwSnaPjGtvwWz0tCeKwfkoF6bN6NzuECbpBrlagv
PTMlFemEctkKEgy/i9x9HpnrSKQFggMUNuRNQhbj+HURv5jLv39NPUifaGQuqpgC
zYmfNeIbeTuh6EWNpJC2joMoQ4Nenp7mA8/CbdSvMw52pHXxg4qkQeT94rFxF/Pa
S7se4CvXmCj+HhiHv86RXmY7juBMaFM0qypvAzl0AjU/yTxbdExxNJHb7CJ2qMHJ
alBY7wlxA5BreL13WqJNH/mFiXr+kX5iw38gMwLv1aBeHXHVkeHqz4OKB1R7ZCUt
Ow+KMLAc1yT5MohhKseQPuu/9z8121ALNNO6lcz8J/41qFfbxhTAWO0WLg1ECtz7
nfw+buvRgu6L7HEeqVlu/b4oH0cvztvA65GBY9FyFIhd6eiBKT5hEHbWj6L0SOVC
ui5KlikBI3nlPrf3HR4xnxTs8KnnxqqlW+Im+Fw3QznABUCfwJMbsAiuZiAp4mpk
QFHB3H0vziqBLg4T5s8yBpWtWJX8oeTojJ1pn2Ty0R58UG4xsvig7l22uB9PosjK
gNVvtcl55+DTCvJSheMTZ2O1ZeQSsKesJt8BB0FmZELHp8hUqzk6lufo/9TtwGI1
tMJ61XGBkwhlfEB5dnx21nbGmwvXm1YxooxOx+MfM6u1o1EvRBYRRBLUXviH4r8L
zRNBe4gcfn2/clS7y94YvUTHIjX4t5u1UUaT9e8CKINSPgdhTwBh2t17e0VGiUmP
l1HwSlivBhGJhgoMqymHG6reKeCgfGfyj1ltIjygMSqufSaIEGdrPAPcpxKtZLHe
5fRPRt7mNzhyLRI075o1kR/dRMqKpQQ6hZ6DOWVy4tg2+Uo3IpyG9LkzAHn5WKDK
g1G4C4qjq9AAqNaMowTDCZGLv66oLJPsDevQyuURvoJFQNoEkML19GfhqTouAkOi
+MFtFecWyWhReBU8Usx0d+K6CQ1wC6nrDeADAxAuN63TFuPcsJ7VGMR/lgIYItIs
p/AZswDnVSyteQGq2revyN6Z+JpdRzihRJnUQ1+7VWp3ND9J6sgZ7MwGsL9+mXYH
E2cjvbbVd3muXan58he/8bRMg3TbxkSMl7pbZqYAK90q4wuC7BDZyCyj8U+FhRtQ
5BmOvViZAencX+N8lIPAYPfPLSVMEaGouTs1ZXraYv0XUKeMxZGvoEDN2O+fsdX5
SVI1yxiOJIT6usJhbr5qYgdW5o/LyZAMqKAtOmRjXZkyPEafbzpmGqN4QBZv10aH
43YWTNeCVj0un9N32UdzOjA/AXWrphrw9FIn2EjDkSqM9jTuKF4kHWblfWkfH+/z
xIbW2XdUQbult3ozgxonmmM0V/H231NNQ4S9v9+Z+Hv8dswzyal8sfKY0tGVfI3q
sxXV95Mb6zAGQ+1pF7sJtonwrhrrOLbiNSaPUHOwGFGL6TiCfIFoLce3XtojBfgb
QinhLJnjpNU5D8QZZzjB/IFTlyjGlDMp9yOVbmfmHAuJau8BnlvWO1VJ/7hT6GOb
Gb4fqhWRoBaPnm1x/w6al6Uuq3ZLtO/exR4CnzeA/GlkD68K35eLj2/ASHlsI2c6
oRsuBgKN28jqG321xvBe8jgbLf3J8YpAakqHabybOwIHxZQBnsuVTB23zvFcoiby
JgYWCMEC1fWx9TgWkpV+fc8n8+qSc8wzcvTr8+JvyaQNawB4W7wDjBGdt4i3nmAT
YCzlCa/sdGbVAjAluRCaj+0QKPw4fJF+BSi2Fyi2VsXI/qA6K9vs9zl9hdqe8LaW
Nq8mwxfUEfuruDc5evGlTceQ6RprPwahw3HlNe0yD54eiLXjfLxdafb1gpXRrH6w
q1GF5QfOzR0XQVvgDQ7h19OczDAqR27v2m0m7v0xuBAwc3hoF9arQKn9TlDD0V0T
gH0kg+QXEwfd2d8IuMYsBJmTz923iwU+dAzI9KF8xX94jCTyAY/Nfx4Y4juIH1he
YIGzK2OYMu5K5bP/PqEzcJTRWcvUT/ym45ee/j/8acgzq8dBcaiI+L+oOB5XMjIF
JtNFCMG88Qn4R+tY8PFsuiJlaXQTSJm9oPE/UJ1vWK5gfMSa4lmUKzWvTENI9SGv
d8otPAkJOmB8LeR/tcxJu5Mu8/U/iUiMHTul351l+Zx/1ctuT8o3Z7Q80s1x5ok2
vlcmWic2ri77k/vw6K5rmxVn8C/SChEg4NCitoKO5zUxIYcEhsM1SW9EbmBdt3fm
KgjG/6dS/Cre3qfyk7XcNiuZugp8wF5A7jZTcTi+AYGw3xXaG6s4YjJd5h9QxGj3
ELLvdmBho/Pm215K98Y9/M/8UnYcANErbwNXpRj+uBqHIn+wzEDOjHg35CpjHNGO
QnHNwP7ht4iDTo4OW+8M/Rr+Jl7aDcuJmbNqi/WvWQvzb0Q5TS+vy5sNwOKpB/MW
EkUP4FoEx0K7TqPtgNEX8xU+7Nx7lDmVxGV7G0ZXMijATeFtDSUI+3H2cBcSH7vy
IDWp/pUA6jcMW3Vj9VTnJF/piwoihnzuWV+MS225F83zYVaNFoVyqdRJXBRbNjV+
zLA3vjoDMNSHsLWhpobw8tvTmQclxsODMjyUm7N/grmaST3KCFeaAyBvD07DZfch
L/vqF/w9FfHZ/6E0Tos/4InEpWZKbxiKnV/5BeBWbfcKuOj2VQ5DiZ9PcsIjYo44
Q/xHJpOIy5RaimAmI40zADshfUitIh0Ryzt5m+DyJ8s9OHO0RQhcWuCWMsOlu4Vy
p1OlpgfmaL63ieevRvozKQSk935a/XTSTKSZ02OFNwXH9iibfqswyIMxHUO5YRcU
JpVhoHdzfR0Hd1UfbDT/4bPOj5QSCrwqqMLPIULjQzDKrwGs/YMwcPL3ArNp46L+
ESgKGQ5/pQF1ouRS3Mj2OPHNiDkTL/wQsyGaGx9B08AwRFaE5JwN2CEAN/NnAKKG
810QCBMieLVNdsl2ThLqxwAH6AZ2blWgE+FdkWKVHa3dFU1rz+0dqXhI2SkL7IZb
raOSthEQnymRlHAwkmALxMQrY6dVmBzjI4jd6klkdNHYeG44fC2ZqFmsCTH8Aef0
BvXu6h/ZTyhXvOnJ1JeQuWar0df9lTn6N6raaX7X2hztQ83YgvsPqajOB5purI+r
Hx6CG8BPsKfTVLMBwJ054Ek2gWn5Ey/N3bCj5i3kTD5oEMorBPC1FTQ/DtscB8bm
0LtHxdJYWH1KlNwRi0dD9xjkDZ+/E3cyL0eNCc3I9rGF54k2vghE8WkajeppdEM/
OHhDgUc28/NGCldxA74SUkQBr260afQau8V4miF0tBacsYtCggTn7W5jm0QxsL/w
ZsdqgMPj83QMRsaHDali0ktn4kk1xyZVe+MXV3jPcQsqBVK3DT5JTSYhFloIk/V2
RpawDg+yHQlb0sAbVetxDoh6XQG+r2eSVrpSsSYtCrQsdKMicV2Ya4OyWaZOAodz
kaSkg/1rUK3/uA8RdUULP7jCiSRfmiYISmkdWjcKZ9vMEH5PsBckPf7gmx2Pk47V
LFtTMpyeXtSVXQk/o7X4SFHyIr9efND1LU5HqeNzHXM+acJtd/brESL4YqD53izX
Ogz2/AHZ3vUZCAaZacDrB3VFCJFBykOHSI4WGHqbPngxYDqQnYPo1NLDlEAK2LUM
m4BSkd7lAFHmb+8S0oQY28glMVz/IaeJu2YHuQMC0b50ZPlG9awc8HSdb1tppd6D
pNNO6AkzVrrsJZudOgkRcUBH+GPTzc3RvcfeblZaar7LdkmUmQ9Vh9ajTLUqaFDk
5lTmfTg3kht1A1AIrpfcoJKIpAbuJNzPAL5kWayIvrlECJlqCTYf4lbc5qZK1c1p
NnMBRXDDQMWvewpJNKQii8ngCpRmjJc26WBKl/nqCWznIhboWIdeAPzbwSbCFeWj
jNuVteNtsRwmWPbAUoPE/IXcrMxCSEPbx1oy7lyajXZ+aNwyaqdFu5ZhP/NhJixK
KC9Idt6erCVqy+/Q7ZGxyttBPBpQt7mtNVsMgJFVLebkXNyRUpZPo2kpkiAA+ARy
/FqtovAekOiYtD3TNEb99SShIblE766jlC8qrRJRKx44wnAWMyIzR2CPZDVgyf1j
idArBN2S3Vl5FBNrhV+8SOG5WygqKPwelq5TH0zpJEZIDzQ5f5z1O/M/hD2+C7eK
cNh+BkleQOd7BajrkWsqcpniLocTzkLEZQ2HPLH0rE8MMgwsGA2iW5QF3OL4LsDH
neInZvGwLpQq9qN80Two9NENGusLvEWAW6M05qf4pYZh8rzf0+fGDdwPrnoUxswZ
9DYEHhnEBdnLW8gFE8H9gOMSMvclJ9drcsxUt7aR0U6mdX/OuR8jBeQI2LeAbC6P
dXk7aEbgxFFiYMvQxiYvc6VkRBNxzO8lfAnrv6dy6eOLtSWLTPioXMsv8fOZ2v29
x2hASolvLeMS5WABmBeq9kemeLiOA/geX3+aGEFJQfXtCHH3yYAdM8sAIxbnQ3fb
3LFPCuPiYbfVvik0ZxnWQI39ICGEmMvYkXt5qxP0m2sM1oaxRcC6FE8yprJNwQXx
ttWyrlJkR9YCINEOpO0c+pflEjQwggPWd6VPtsIiDUmngFpGUrUnPdWrSxhSN7jm
MoH5Z9w+tW79qPjqHGnWAa+FRjXYygS+rzfcX5cStku4o0AW1Clc5OTq/vMOw4kV
FmR8rzv4X7CxLFM4fQlC7lzKoaf7UDi5gckCHj13UxqbV9jfrarBddwZPi6hlxwJ
dl0JT+HAJXxBSINnMHu1utJSjCHzrLIn8ncqF+ZeEoz2J3fjoW6eXtDtkFNNY7TM
mqKKoWePJ2rtjJ+WsuquF3LPrjTyIU4wSIIkt10amW2wcHAiR4g8+xizgE6sJ7g7
ZL52+bpEdOL1itFHRvekaFRPRFolapfQxP12bDp5U2ZBhthLxhDz4FE3uEH1ev/D
e1mP2eskKopiDVk77XmQ8Jm/Uiz7mwewRghZrRf/qioHoOV3pY8pJzGtgXXbe93t
Fg1cuukfryXiPbY0Y2bZo/v+TGyhQPkqaM7NUdjAqQpItP3rR5//xEhpY6hlztJe
i4BCAssfl16xN9BvU/O/q5QZAoh6meL3NHvljB5OiZkUYtrimXD4CDV/EMV8U8H+
jJ4a1WffFyAKjvhZlTJXxClky+zU0kAeJ2gdEwpLK4HrMWBdnKtigeD3OEDhzj33
h2VXLHJz2ciQim1IycJy11k1R8KCZH+DDwaJrjKyx0YCyu3UCispV98x3fDKSwkv
ChpAODFjJAhSsy9k0qiJs8Cvwi4NPobBJLVTTM0IEc5iZUbZG8NNRSkPUvfzM17b
H2oKGDlJ4Y/D6REISw8zoqJuLd7PYc2aBtt+KhWjyS7n3l1265A+S2TOKlrLnJ7P
flHQ3B8za0NOynblS4pZZXJg7xZU5776k5/5ZfgNfUdAe3NGiTuEyMZxR8Q1q5XY
/ww0ZPYivkDTWs1GdRWUW6fyO1iGGe/CIvNthJWDd3j2BFKUtKDZ58xf6WADsrI9
wsgi+luq/INj07XSHaRRg5iX17Z2g2+7M+fRWRd8rYMHUsOrDURp4S7PlF3RLrbw
GgVYXPlLJV1KkMYzFnj5w2knj59bsB1U+Q+ujkoOsOxzuqV8UjL+3ai+O0iU3QmD
D2CND5BqaIoAHOdcKimnxFrFErKcLsliFRrPeJsdvl7Aa4qBUF2kAzhlSNAdD74O
dBI41LWZ6gEClu7bMhUXi+9XpTAEPWlAutiZV9c1CnAIPC6uH3bgcKC3QnNzv2CO
TWhHrlN2gUTHhJjdFaDmSg4wA3YXjoohvkiO/kjqgDJDSjkiAK6Zb3dLjmh8wdNj
b+kZaPXarDND/AygsjuYj/pUr29pfBtXoWVeOlGKhW/s4x6rcmUTV6ESvp3i8Bex
dPJ3iEl/C8aHqxUVTZjffEDJwLX/L9r1ez88SDd3H0kXXg42WYFxF8fwuegxvKIA
FPCRvBL+fCV1y0XVewmz+p9j9h84LQRUb6cpy0sllcmRzu/Nu27RoHi/kIn4zyfV
jy02h5XKYu2P4dDSUOApTxqW2UAhmEdA+gQkRTwSXq9za0eqQE/Jkmxv2PEkwtmM
WMDbw7z3CK/S7ilUawqZstZk9DXC8AMqGxGH9capQ9zgtxDICYApMmDi7/S6mkv/
RhU+hBc5ju+NGuAnHN499rd9O2XW1Y8ZeCKpOIsttJlzSq1+kMz9e62ZnOH/OZ1y
+Tw2Fn7aUOQI0F0h6cMPXQ5SJv3fI/TIJlcKCpM8saqNW10MK0HDIMHC7/5/aMnv
kALdEj3QQx0y2KgWrSqpPb5Z6EVZDDOr3cGT1IxSWQNDtmdmXer9c6Y+5+8OhwGu
MclWvgZ1M1athFoRYmGXUlYLnK3w5QGyna22R9AuFXl69NFkLcsP0jJyC2bsjbcw
+bB9aahd8jhnl22jGGEqghLedO49zdI0jXghgvIVg1IDJ/J81TFHu0YpHj4Hjrx8
qx8lcHglqlpq6dJq60iI9hZR7NPb9nVc0HrLvUNGH/yv+bBuggEgGiTmlx4i/0wI
NCU269e6Ufr6NkhXcZeW+qmXamZrZNpy0QJkaFjY3yaN5v0WdxCgRE2vfkNAI1MG
cru6XlwHCpTBpBDW7emxK/yTshpWHwditFkRUN+odXKxVcfdPWv1ftykbo1WsFlz
TqKa2bXWOX34QAWhMG7QpR6v1BgJ3eRsku/G2VgrTGM90/d1MqjkFPLOYfQF99n1
1AWFQWcraZCRVgqOvwxICGMMxWVyurX+nbi5YJZxAqsDonUjLLzyePEAoOQtZLUM
XUQo4sRUfKSSvAaMpnq8roSjnTR7lzGRnlJ4KAs/l72RDerlONrDfS49o8jqsBAF
tl4qt+rYsIGyooOtMROclkmpfpDBGV5d5OKOUlubcbCkK1TRzysjcBtHGruF5tP6
1VGOt0Dara7SCbYYXYNciOoZkbGl8kp45W67W2klbSefdF7PwPR8Fy7+bpkXyoRK
rzNSFofkFR62sfT+i8j7cMe6wm2Mrvrzcp9qbfjzbaysAxEZPzDfEntMCTv3KY8A
vOeRguFp3o+NPlEDUowPGUUQ5kCx7Zf/kIYD2d4iOHoYoRfoypI9Y1x/HV+cGS2I
KusuY/961e+1/rHxaposEGbAd9AmNwzeYM0PRVv6tVlbe/wwmHc+F8Im5NDMc4Gl
FY3g19OP6gGPJtmgT2AxvOpxWC/7RI1+lDLU0L4TTJ1PvzAWD5cSN0MvF7ckZKR6
d2zFjFqS+XwQXdFLbiSQ5fOAk7BMWjwV2ecpve5IFHPNJSWQn8ksOeddRBmDG9eC
jjAldTFjzB+HTfzSM5f+neNWnotwLccT72Vq60lJWgEWoYsS/WwxsufzVaCMWa9u
qIM6UUUJ+e7pF278i+Kpw5oxf9eGlWkNeQ0HYmMgxvOJVjd8sDMWkmgh/7kd4c7L
YFpZO2YTPTmBkR+3pAF3NMQfDgeMffJa4CqHyFN6jD3jS4R6RZ/0+ErtMnMvIE2F
hH71prj8XbkGHCtS8d+OmTC2+aT6DPodL70G2dFc4Xe1Kndn+fLaRT9f/E0RC284
Ab54C15N+71e+tN8okKn3/UIi4z35rpTrD6Ubne/lS8AMGW+AK1dvVGxPrWWyuEt
wafj7qIYqXqVMDsao9j2tcoxE26oHfHSM3Ih7r1ksCImDy+WwpyF9AmfDnJi57N7
jaW5zSal/13rOkQeWgKcE5WiOiX9NjhUSx8T9VR6hEBxj+AKmKxoeeOIo7hW+G6b
KOgLPlRAW836GXvdA4jjuS0cYzGM1NdhDJgXiRJVi/hOXwt0+0wUqiWIBngKN8HV
D9Pjwrj8JeaaCCQdUjl7XYVTMlIFjquudq1adCElHOg6HfRSndRQnEE/2GcQuRWc
fr1JfOPm3VIHc/IcK7ek5Ku2WiErD5Fvn4R3FfyUpCOCL7vuhWsw9qPI9s585JPq
iS3Cl7ekpsLwp26masaXkswbpfBvX0odISnhhkgKfXKfTB/EdNJ9szv17Pwnj+sG
BHEKW+jp+vl4N2Z2Kh2XT+CrhNyDheZEcHUBV1yEefgo81YPzSetwpfLZu7oYlHS
Uyp/3Ht+RXjc5KQvoYDV7rdkSmjg1DoxZkwBVcqlD88po1J55sd3grphwpGjB/0F
+8hC+c1WlM3svPyvyOYpRlJHAHXxdaXcjFO8Xc1gF6imiB70v3EueVI/2Qz6htmW
Q6R++BuuP4JC+5LoNdWRPQ7QZcM4J7pub8wkILMpaCK2zJtfB3cM8e6HSh2zNm54
ef4ORASRafjjggpfNDpxWWBx0A7MXUNcencr4mEiO8VYo23YlZfoVdKZ2l7futB9
E+L1xaNZdZKlEsBQQYql9v3A1K9IvLNOD/RYt7E/mB9lZrBCtMzTcu522m+/45vl
D6QWnuvqLlQ+BRgkvktWOG39GQ87DJ2Qp7CYZxpbKfKjsvh/bgtZvbP9wRG1hCJy
TOUZDi2J+NBdGIAbuvhuEl1yW7VxN9kWdH3eo4wdhgm+QLC5Th+Q3RTzAroIY1zE
ceuTWJKS1slSBKF1vMuui7HKL8EQo33WyU5P4EDJaZvmNDhl3yTAVooLhbFO/o44
0+KoRLOla4oCHvb/eiBkVZTOKSKMR29YLhGL6RdB9jk/lY9D9FoQN7gEPQLGiDd2
QAyor5xOfZVKDIxRMbZqG7eOzVZrSPenk6FytM/QLk3lJrlA/JwTddWbzsj7I0Al
/wGk8sBl9GZkkOBKguZNGN/MrAd51VEDWm2O7IvuxcH8h9IcRr5i7CiaTm9mv/vT
C/gt+rapbNW3lVnm/e8+3ufl0cscoTH0T23LKjs/jj05IZ85PpgzXyxDNtJuKLkD
xEGhGf4133YbkIzJZq14lY5pp7e72f4UXMa4knbSEjVo1JrlJ2d/gS9O/BeMXu7J
/rXka24DL1vl3r2drdWWASZHDNa80796oOIAjkpRiX0CLNbdUAHYJCjDzp3pn94s
vjyqkrT63YAG3oRxQae0vL9twPU/Fh7ISNXUrOyMPrwO4J0kGu1CZMI0zG98KjSC
FywIiLTBzm1P6WWy3/e8UxnAigp8shHB2C8+MUBTyc4yUzlBmaanDHQnSjQ96MQ8
wIH5k+wmvoSk8bZL9YpFvyg/N4w3va3Se8OLoQZJua4hFWo3PDjzSYURQ38J13Bi
SsJ02+jhyC4wbRP+ncczGirCZkWekhjtnWuXx6cYxioMlrbr8CRThKMJHqiDiIm5
mPHEZ8knMDkLFjKaTZMHQmJr5XFzCyTeaJopZY5hyDEFwpWJw7hU9zKEy/WivMJI
s410mdOQpntkWzEYE78wR8XVv4Du33mGy67Iy/G/BT4kbJrxTUxcm2gTOEXGwQJk
4V6gBw4VMp3Dtn78iAMrx2m5SCMppi7GmQ1f2d2TTTuQgWHL0LLfs4qEo8ASbtLO
1PktrWzsam/XQnOi9QFk4RFX69szLLkqnia7IrseTosHJsh0QXhFNb8pbV34areT
tpH27POnXeOhoL/JOJngDgAl5prk+OjUTGjGUnUC6DkH1XFoxiuFaz8rwlotTZpL
mKHWM6sJQqCbW8aGQfFdPQKd1NbRQQRLO9VvpahmRxt7Dy1ygwSoDPk6261+kH05
dcXDkiYt60Y5qP7v5LCWrpk5CbL2+f/T/jW8uHeGX7RlZTzfWO3R1My/Nu7kjpx0
Q72G6qKARTyak8G3E/vo4U7wtfTGZD0JIQ8EnUmtXo3cKyy2jUOTNNltIELWFO61
Ct3Kss14syvEC7bMh0KWvz2TGVReQMoHsiAneC3cEJR2CsgXx1ien5RULl7h97N7
swDUsa5+GKOIw4X/vbOCkkusUFI00bSIZmHXQMzXDZ25Kuz48n7KFO4E2JyrRwZd
3rFkYtOVngm+6fc1WZiKEZjULgrgXxmoFA2saw0YuhXts5Gi0GTeHR0HJr3qGmkq
r3qzDYIwJa/7L5G9L9dpucMH6mAk2fMKOhZDA+OSZ7Aaud4AJpkqKhKTy6eRaVh2
vqNGTmNll3QIjYuqA0MgLeIJ6tB/yrAqx/3N656tzNcaVPF+GvL8yV+o8GZzyR+k
qx2LCqG4/Y147l6hkwIQaKIPrnI4UIa3uj0yKKkXlNnBOLLzsLs4w8n95LT60ooK
PrlnnMRH/kBOF3UADGe8a7ezFvZkwqsXhj8HXdTfPL8rpdDJ8MXBxkcU/Qoa1c18
3SaBWyUhSeQ+tYhUM/l2PqBHExrL/8dvCR2R5RjqeV3FOpHpMaJxLirXJtsz/os3
OR1lRc51iED18U5mu+HTLgLt1V3+5pKhetzpA54w4FherKcsjIFeBI3ji8tLmpIs
7tO20hmtD5GDv8XANXVgad/3U02zIhdGH+oDsguGcnlGkdoIJbyhOTAl+s+pdDU7
8pXL1uQ4hVpCJVFjoeeaQ04ZxfeNmTASDDrNVtZUGNnnLajKV6acTf3SEvyOSZlW
a16/OiVKdWPbB+oOqkvKkvuzbQnXvUsbF26aR27/aif2J6Xi1IDHVJ7RPDrLODhf
q4ynfKtl3jmWc8M8TnTb4nevleXQM2IFLH/XJTQn+tDWD7260uhW8D8yx7fJiLKT
Bew4lO5a0aPVIo/wOlVM5bParP9dgX4Q5ZwSda4xetq1HuOcgvkkhIO2Bd8u+w/K
+cveAXEY7cxDylKiGbFXcIhTw2bzDECwaAM924MB/E/GaesO94tHk3YzfIlsQfA1
M1Mau3VklLkXuoJoOV1C43ZqKSZAbmLlKPNPGZfo3fHkVEoMd9xf/YpAr1A/C7WW
6fzN1Nc+vuxqx7JmlZvkUYhv9dsI96A3nY6/VicALhA/+Lhk1VyjjQLRc8noTNSz
bQCfAloMux78pFNjUiyb27WgwWtksa5kHWBH7uqemfpKPudrPbyeDacaj5pzoMtj
Ja0zKhUQivr51GZLLLwuJX5SDlaR5pC+IFOidYMPWlxN/SfjHeNoaf1urnrwAuAi
1AGbfbQhM/6dnpGgys8hMDkcyogvR+LkdF2f7ZWBAi39Sc+t44ydz+uj7cRadm+U
U+2ADwMf56hcpH91SRhNdZo/z/h8MTwXOQYuSmzBG8Uu+fSmGDBv/vXGcfMSNW+8
Lce1sZ0/y5rW4iw+RS+aE/jrsxsCCqH87/XiTKSSTCTKVoEQaW29spaIbPXedqVU
ydsPSa3DlGUEe9aZWT88wADhyr6aXeiacAWtKmH8YizVD5pgLlemALTtBQcXMrr2
LCMG1pP3dCX4viIWw7ap11g2aqtRXFXxV+5BAX9cypbGCMDDxXYdoZMoDUso6xez
nOKVsW2nOe4sBkfz9nNAHYECz4dbqgk8up7r/vyUp1OjznbltXneYihmlmYC9c1t
AtEwP0zbtqEnv0kfv+iGlWQRS35gvMoBnGe2Jb/eD4KnP6fJUbsPCrkT2/b+lVh7
ke2LTBW7HYDbxWtBXbaqWE8f90uDT8FlI+A2uWNnC99WhADNFwMFYwWmL/gz0kuf
hD7wjMJLZfZOGZoTMhU5TUFDrMAW2ejTtMrCKCMZtyUSaFfOl2Yr5ugo1ctl1j50
XC/0yeBCkYsEpyL2416Jt2iFzXtTXrQ9B777fXJtEIvPumapL2Rwil6z2mdP7kAJ
/OFcdyJyYClBYnYUJ7VpeLns2AF2LWa5UulfUzhUQwRE5opsZK1QXH1FbXJzZWyA
6yiAXb9AVRiS02Lcm3byyoBKvBQlXlMipbB2uTebvyLZbYPB5oIZ5r1f+vfcCWNs
gx6tbuSy974OtzkhERLqyDfmqB98I/YjAnQDxAUlC6hElmdu/VTkk+XB83wAVrHo
gf9zosnLtxVJNrdMLL+O6910AcwetsfV5fDOIxluMYuwbuCFS/FwJPIcWeGAiQzU
BOrEn5n1qKlPGcncr50w1xPmdare8dEXi7AgOicINNDAXwtPpYNFy4Ei6uSuwCaP
YMMYYut7tswZk7VpSaQmPqPnW6N3STaARLteGCeGHCzwnpQcWoIR3SIY2nndigTZ
X9z/tVWrzn+deFGwsA961Hf1Zjyhmg5jC3kBgbgdsomfAm6IGySju5skfYf1nq+r
UbFzPRPwnXmlSLfGvS8DGSpj2En6RzjPnMptgMsk46knXRgghxAq7muYc1F445fg
R7tj1q8YuRPMwRvLtGitybBt6RIFD1qxFG8PgTFppKSEd47CmQkdJyFvntjgoz8y
jLzXvj3q1L0s6QbNuTmvfq3rOwOSCMh+HnE0gVLVmyHFn7R/UY55FeJJUa8f9Obc
T+iMpsfLn/6PrpYAZ+e6NqsnRrqdwUVNrSv2JTC1JOsDo7Afo7w8W2zmcUMkvqgo
3AsSCkg2dwioHS1VoUOyDuihj0mpdfoNKuFply87+oq5W/7qJj4T2FvYNwTroJoe
sBPjA86zBvi7XWm0Yl2zH1n6uIYShZiw9YcvuosSCiYI9CwNbmjOjhDRrwVpQTHA
VcmmG8QvBYfRR9HNdydVwudUW8f82L7aiOI+jS+jCKrEJdj+Y87kgal41nm/ZjmK
mTR/4+UF61X0QzCVStQ+eWDsvLn/e44tJR9KD3rdus6JLIyq1R/3ZmeUArgLY1J/
t7FHREFQxqBvnWC6dhORXCMqX8Ve9pwrVrpQfhUImhgt7QHgL8cVXVKNAHeImNs0
ufSdZXMoK29ow44ets7Z1xxp3pAlTglPE1lskiI+EYXHnECX2BVnhHXDSSB+j/wv
QPedhDPg4On6mnfDR6XD1OxE/0PyHiN2iFb4xzzvQPv6z6nVQUoKmN6Slvt8zguY
PjVc3F1zgt5rrnuVSTnITaT0FqibjwrQO2qKPfYkqgY38+79z966bl6JWtxkbRoD
5sKRH4XuRXBjFpO/G8FdNW4Hg6CAsMH+ivX6mJdxzmvtu0JQQS02k0gyO5O+6iG+
i1tTjP0L6jQrCVMgJXSSQwgFNByMptTssnT8B5ydAbc4vFdwqejgoMLVmUT79UkW
4VUh+qGPjeoMpuLgdZsVhNMfaLDMIBMpdAbOWz9oejvKdOazLT06sHL0EEF4XQOt
ljz1XESshnEKfxS3QTltAik1Oj9c2YP1O0180V+yvYFDlQ8k/E3OoPpXzGN2CG+f
H3olbqHxNAW+63XTC+InaYOo9vprTPYBIEqdEQ3feoGwDJyPy2rb607sfyUUAJWG
tRcujQBz/g47Fm7kIxu+w8BZTnalxCoOKmZtzJHNK+F9jkSx4Y5dlm3oC+mZZvKh
RXLmD4O0gJgQbCDE5+WfsdBarsUgfeTBiK5EHDp1/B2rbz7RYF3OFtl3HEoyaONr
AyGtW05LRwvOR+/6ZdQZ6D2hxtEJR5nA3+xzoxb8OtVwuugJhmbqic2O+gTa9zKm
hQWi1f2EwRDHPQUxWVQ0j6GJmeTM/MrYamds49EN4ouviOoG0Cp8c0AtjpZFdfc4
QNoOFdAEmr2cX5oMjBUgK/vPjKnq4mv7px7cVuHLBZszG9odGuVnTgxZCy2yTJPk
I13gydT/IIC0MusG0oWw3Qjv7TmwR43i0daxv1c3Yiz+iY13FDLqv8CovsAYSA0r
p7nYIRLgSzijfriUaIexvwUA98zg/J7yoB7m18yk67WqtMEv3RFRV4Zmpo5UxtM7
k04KWEpAuxNkJLFbMdVo+WwUF3npUQCTZl+c/j9JSm/WWtwYzzh1mqNb+YnOMyXj
EJTAQTBzmFSWBlSrYKRQCyeVDdw4oTeFw8DeaLcAq5pffsz946o68IPrwr6XybEM
wNhiXaQuiAB9wciNIYKvbXRB5kr1kR8OmxRONzwSEQOHiq9JddHGIRr8ZQQtGcNF
3DPgQJ8QVYn/oBJQ9zkfK1MA76VXOXgcONI2DPB8TiZqLikRZ7qPE/XlXxncvcBy
SYumaVo4YEDRos+OVayqSTLoyICSlJPjSVa8dIh9kCpxQXMjDGIqUULDLCT/+fWt
IoM/9NWTeAtQaYaspNdppu9nqIyvfa9focRZB2YTvD4qA8rzJDjohoK+htqVwfbs
Unka/XmWvLJwrhA8feV1Ea/HW2RN4MZ0DMbAlUIRwJf906D5ALt4smGvNFghOTtT
D+ZVK93GaMnNDZu3C40JATkWmDbj7XDTbpHca72QT24ZEEP+flb/Mw0VarHVy7yc
eTAtD97WLA/q7JqRCqzTW6AYktncg/GqW8CktrtqSIQmanz2N/ensiI9u7HmeSp4
oiYQMKV1kanWoPFc3TQzbRCDAl167a+w9afjE9gGxkfz2X/AS2vfLBrdKjtmi9vV
M07cyaqeSv8qq8XBjopkxNzfsu/BVZZF5ZJMC3QRFkD7QSEXW9PpCzAZM6gmD8nt
peTOvA6/6UWWISuqtdl6AUUXffFklt/0rJT+ARfKYBZhZvVmRGKcMvd/5QhCQtfs
iHB9y+eUkkMAClieX3KDL3qTPQ0IDfpEBGSZGIFjE65hOmC9Z5/CM6MrEEky/d3L
m+SrQmOXsVesc58XUdkJ8tGMneM9JmHY3R0EEkaU1Ktr/sOj2NnN4ieuXdAS8lJT
NWyZ/72V09ZfhJYO0PAk3Ex2sL0EU/UtcoeQrwU4naKjhQT5rnvsefpyMam2z6Tp
552aLMgUx3KFFal/aYkpeTQjX2s8WsK9Sk82ksXAeekmw2UYnwIXxhg3O1HxD6hd
WbnbB69+pj5QH2Nupgtj3dBKIT5mWgKFsBO6masiUrz3AL3P2/bNbCdK1tnTzPMH
6GHzthXACeOE5oQlbtYD9wgUsIVKC8vmpF0GYNOIYLtsEBX7XDcxwUAaYJPwOiSX
hu4ImwjpmfjJty6PVzPk12rTogvmINiF5adkdfvin2G2uHHAbkyLFESVPokXVIYE
Lyioh5n8taq6r/QwJbcld0KUcoLDOIgnzW9xT4ebsIN2RS4C+HGfKo5dmEZRgeMA
c3fWhXNzvAFn/snsfaVoM1cMaFhLpBZRUucUdMh9qaLwYlSa/HX/dt1JqELR0Ja6
6E+t4NKUX2nlBnn6WMaeQKglUFmn0zLy+Bz5Q9zJ91BvFBvw6OMl/A3yD4/P4TcQ
vXD3rbeWIy+6YEkdAM9LO7bdrk/iOupXsogqia7+mZqv37wbeR+d0FhPQazB8bXb
fV7zSHM+gW7eeXQ7wVMn36Gy1W4m1Aqkfa3hHgVsaXRGKxcEN9+R7PKB5d/o/EQj
SuAkj7V7CxcmBIf7zhwGck4vD/xqkWHztiyHKRpRBFZpXa5rhgWCdDUdgOzclg4U
u0UYn7KqSV14pRkK6LFANXdaI4d5bCfBxDjXkx49euf0CYNbDQbfdYvGzc3VbTJx
sKY43TJyF5kbyy+9aeonLeFQCwiEGWVJarDJwbTO4Papl8ZOXV84dGiu/cmotiGK
23ODcsRGBZII077GlfG4Kz+QlSJ+wJ3u+JKDRWeV6H/5W3mViT3uqBu53q2BCZa9
TNJH/p6yDn5fTlm5BFwhlJ6zPVO9CVn1SZsQwnH+egpKX7lAgw9anppBLQe/MmI7
Vg/B80k3XOc79pxsvnp7JRx0uQJf7pf7fJla7MYi7XrBkiYwuNDefZUwBpJXs6SO
Ul/BxQSMH/Ci3wSz4yKup6wms03GvSXxonP/VOV2NVH+C2PCIBCsLpFx3XpKvUp/
WJDKOq0uF3zW8xuwc93mLBY87I3+9qfzOG1HeDjbPxHTvg+LXeG9tm/k5Ae+FCqI
AVJ7iF1Eps7VZNkH5jXKLQdjNK2tSry5fyc4cLW5nKxG0no0zERbc1i5ePe6WZYm
WPgQE8MESoKRvG/MGsH1+Wt/H6W5XXwX2s4s9RtEeyLUyjcKUXHcgva7RcADSq66
VPt2hTsYp9H5BacfMvYbeTV/A3jAKiWmcIFjgS1JgPbF8LzljWO638mR0gCS7c5G
trYln3e9j1iW4pK00l953xApJ3huy4kRvtI9ujaR/Kkbc8aa5kUiMWvlWQad1rgR
d858B4qK1uCAyD1vWzfY+yFgAWs8Fw+MMky2snHFwZyrpptccTut3DiKQgnMhUxe
wRE5A0ltTDfSwcPEf0zbJQi+/A3+y0WH1GH0/HhgIVtk01TrRypHpDtl/9rupppA
eRjCkYjX/04HAuJyMqNO3U01TWLJgPvjgKdj5QDPNrF80fM8o1OEQu93RwxeJ0WL
Bpyv5+qia80oyocDTWzqA5cysUHNmwEPDDwUsEblGxRb1OAU2TFE+UWTXIAOQ4kX
z3zU2ytAU81fBnV61UCo7JOwVqysq2AD5SQOuEOfWWgxT93f2ZcH7rmloQKA9UXH
0pLqukXTNhkKhe55QYV/EwsDVHMTU4oRx7/qKXd8csnMrcmJYBqv8SUxbUj+omyg
stT77XbFNIlSqZrTD5WP4fYBYxJ3lWf8/Hqzb4q1rMpZpf35wtcmpeYfHg7CtQ0y
pfoKnMPSNPgXptmhMVQr8XdtWQ8CziPWnkSFT3NjEATrn2vaJczOyqsK99aL+hSO
Hnb07UIKxKqbIAnneD6NKiKfRysILiWkqGK+IxiZi+PTnC9gnaogjKaqg+sCHp4c
rgNGU5fuMO0Qc9YvuwT11rUJmqvl7Y3Ui4rFO9/KE+WSLNchxpDSYWobsqmIg8ix
rbb973rj5sBlRahnWToJNAi9C1Irgyoq/Ljm5Oe3ivEJdiEnDbOfoGRcePdxVhds
++e8STi4of+Gv7C8RMWQAgRFJpKc6lmB9J2QqSF95sL0Mq2WnrQvToUaphP87n5n
+hbnNruRkZ3ddSWgzFCy7Eyp6cqzl9zhdi0Zle/OnUeIqvwYWL8WN4oNZwcUbeji
zBrQoz1qVo2q3lzC6n0mIPI2Xfs/X/HnZ5Tm2Eq2dHdHxw73gJE/T1nGWznhNFqQ
T1isBV7FnW2MAcs2qApHE2TF3u4Hh0DLMDSAPrWddgtk8mtGgUV1RR6BShnm/iaF
VXN3j7H4bTtI7rOl/FlyrXuolpS8fFUTBT+g0HZDRK+oetXVy9ibB2L6IjZuGoEl
BrXB4LUq82hAwISeOSbEFVZ5K8ntwRUGRO8NxdPUTNK7w9MV6TtRY5yGUtZ26ue/
pNwHAH+pF5TyBjpGcAtLwHBfdnRoqmuBDBqqMaMTXg3e6tE8I1L0qE7p2ozOB6bv
7ga8AGoQE1C7nFm6hq27a4OF59izTNcdcDut5+FxMuny2y+0QZGbh0/AFN3s5JYW
qY6Sp7lSICTQO3nAi7XJ8PlTvM3IX+X9IqcABbSHRHxZs9Zt245mB6C1/cidwb4c
7H1mx0PA8cUTqB+kCN/NASkxmjb0SiC2AEfl9lqVl5dMpZ2Wf0dGrSPIZiJP32GV
gelaKdfLMLyDNd0UF0pXtcGKVXt2BZnAiEAp4wnP5xM8NV6PE+0OE6Hy1Kfy5HU0
Hi+C4v0v6d+tyUuFvNhm4QonV+HxhWhAoHxNU80Nna86Drr99Fj7Z7bhNMPtgX5w
eMs0LN1pKemTYKak3rzSlXFHZJPEt0d9CgYytYrYsUKcayBb7vUNnvh/NdYlr0zx
T4qw2+B9oHDfWQLk5p3xoY647EsqCX+Y2sNDH/JDBDlE2NYaZPtUqhKV3KDEEd2r
bfOmk/dfUf1mQO2dkdZljell1G4CvBcDzQQM3ksIzaW1hOpnZPMxsth+jB1AoVpT
jPQl7c8CHjmbiSKilYS/BEObdxo/Mc3e9X5EWpofUc2j5tt/5S06YkUgBXoxr4Dq
VwqbSCJfit2OUYvUbTjbYolT2CSZzJIQ/3RPC67mdqy/6x8V8uyzNH+hpiRJxFuI
kfHbsN7bPhAXXsF+C7lh/PdpYkoxh7kGg+cF+a1bDqRZj+CaWDBK9zQ6B7qYl4YS
fk2ktioia8I/9o8+8jP7Wnq9GrSXMsUptpKLQePaQwcf0yBCRSLsJ06p3PeY0Emy
PoZFctUCf15wfnsyqUCz/FZ9r+b8xTMm3VPW7hW+UkboniymuwBU4Bb6W06u4O8D
VrGMvnmU9ss5drbsh5DMh3cJ2zHqwEfmmXj2HmqeC/18GcDB7jImLDtsOTcJKtFT
lTBpoZaIPeZAWaQIGjXgED78TGYDY1qS5gaDWSSrOVDACYJovESI4xtp9EuRxoEX
fgzFh+KpXfQ7wQufTjZOrWHGYOYuVb8gvxRfLaTjnh1GisGkp/01jPv94XJSB3yY
vPJ+iYE7m4T89YfX0VqxcA2xFklqaZFqoKd/JpmVERwLd6YMswzga2kCr00Y+Oz3
Zvbj57jcd1UOrZ6O14XzZQ7roDnPENYLuyAaXxgutwwPxew0RAz2GYKztkGVRNXZ
/+WpDsU4HEexWIxh3MD7i/wc4gwSoqNQNAHDIfT2xiFBa/KbeiLCfWx7LoNheTiz
trdzcby9BvEBlKqfLg+wkqqttgTdp+PELBcLVVB9IRyMLMlJI0jJvHXktwntf/8s
kuFbtOlJh4Yn0H4JDpsuXO0t849m0r8vJZ0gHPvkHa0o2W1TKQ/kBzYFpL67Y5T4
yC2oGeffrReGD8c5EU0tRgfHKOmfBhOPN1RXPnL4fwTp8eBI7q0XSBH25PvBxU5E
+k5s03jbU4e6Ad0NJEbo9/6Y1hKOv4CWRwN1RM5zVGtxbG5FV03DmEBK54Ukpey6
j6bka99o6FZjKq9Fj6RKmHX6p/HwRym4O1H5aXEpITv/4Pc/hKrDYK6jfEdeKSoh
AF6X+Bt9hd7BqCa9HW7kDE1PXP2HqvrFYExuV4pworzWEuXTuN6ojSi0rh1bXm/8
0/yDEUIsvM7t4JuRJHZkoSiYlAGmU/IqyYeUZU2qqsd5HRpLIMhyp0/RgOgqUXt6
YQvwUzgkz/8/rolI3wFroJh3imC6PHm0e/WACzZM1YiIkRiTxWhy/wC3YlADTm2T
oB3ajwCwwc498i7AUFL+xWyrD2oM5uIy1yhsTtPqkOdccv6bQEBbN7LN0xRyqEff
/8lDI+OYuwGK85PtR5fMwH6DYnXfDiZwsSi/cwjTj6qsqdCUMInQPvevgONl+XRh
3cT/XxpLQmiZQWgDuLMAj3x+6tzzbthT8E7nzXuofXnTvHSTHL3Qko/4iTcAM/ZW
j1r1MU6qm5Hf11+L6bKCU6SA7u/2Jhb6/+4WKyP+MhX6747SravegcOTLD46fWPk
0KnUnqQPnRgqo1Bcwy1meOIgHMtIJzHiJeml7fOzAix5R3xA5+TYqFV3aZ6K0rxG
u1XekZhWVcarsAF5TLqfNu/tP5Bi0Ym7BEb/uTh3tqKJ4gQgpriHgJWoN+y7NWwI
X8+1qDXdbp3zXw6j5GtEnUxYicIAleYcRPTjDxud/QLoDh5jtS+6fLyCp2gaGvM6
j+aPTOGoS2WKKn0a3caLg6wT7bPo8fojwZSrsohDkvJ4d38rtrv8eOiCLIcmWYCh
Pe1CVnVQ4Dg7WCZ4+3gfZraUCxBXcgHDg7ZWMj0BITa/nbs6O6G6dOKXZDTE3Lle
suuK+/0Y8tM98hnoAFub7qHpkG5D79dhlhoywMuRQLmr6qmiO2GfQeXhduZ9m3nJ
z/IopmFuIhZX8zveHxoRPN75/cj4uJaAZ3qpN/mXGbpB/oOAXBCDSwEDTOnwUiBb
UPGaHHvPKFr1WQVADmHqNxzNrNGvxkk6Juhyis1ubK0OyGpcx935Ozh5kn6y7ezj
wgZDnl75eHNhxfq0nRzq1BP5SExhuQg0c0bVd3wzZ4V3LH0rBXZYIBStmEYHT3S+
AJUQtb6NprRc2uxnN0fq4F2t3c8sTuKUB7YQ3KOPFPcFPdzgZL0ztD7Ji8vtUCDP
0tUBvBosoEi5kbiyJ8AfrUlTRs6q8CF0AjPRe0yaBI0LBNTbOvl25tWbZPGp1dCF
7Pe0u046j2zMothbarv4X6hlTB+uRUl03Lg9awQ1KhxNz0cT8z8UrOeJigSPvfL6
Fh8Y2mdaIR3cBSmCZE/pljYh75YPhkoDy0pI9mYOlgE95U2kbrZkH9mdNE6S4USO
kvlJSOEBYp4+OOsM+7Le4XWIM4JgNbhw+8sYbfNnxgRdoXzMsqdKJWW9lzZcv7HN
yrc88PYdgmobMkQ0ajbfm0AGiIMhk61wIAQ5QbMYVQLwXMylT96fJmW7hZnphuvK
3tOgrOf9RtKm7PK3FvkDDgC2vKBDLMkQf0k/4Ukl56fk3a1rjpGxzW6TIZ7trJJi
cBKjpfdliY36DoUoGkjkMB2QxTXaR2LVcJVtaU2Zc6KTVH7gJEz0F3VcImdv9vA1
Fy2ijWESBzIbZ9qdaobsQPVVK1l2VSlDBwFqyC3oLxnI/a/hBo1BPV4SIlPAyj0k
7d8INT/9jyQBRs8gz6QXMLs23ZGrT9PZiAf3cecQkbo9p/W0AudcjwCpMd5x8TyT
blyUv8Mi8sf5pF2tYLYm2DU9+t2yWwO7bHFVIIQT0rYjUrx9iWeED5mwVoSADygD
mQtmD7iHZSRw31aESfQ0E/gZl5IEFrUpuIAuYmQc4CwzWCbfx0V70jIJDRA9W+oy
0inCMKZbzn3tG9jnwXe7z1OCWXclE8QGIQtenAnOZ66XA0DgOqJ+hF8LyyKpti9d
2Cqfy84p6VmUV+cTfs9azKP5IgjAsuAarshea9/PrVot18whkQ8TMdKeWkX6kNy9
jhBVRgkWD3ijZ4jCUB64HKQQJ9pEQ6T1ACu7KK4+PFn+CiIJX5FaUHNDG4Yv0HE8
EgtISXIPb+j5EsZvq6EufjD1sT6CbB7JYmlLTIxSeFWy6gWFWMKutxwLgnMJq1D9
04dmmUaCtf3jd19nCL+tlzGcLZViIAX6aC+nW7BdUZ2g5K+yTZ+CaUcs22BSc+aH
uYb5MMuZe0dWd13wWrnzmn+ioE5cKSyjf6D6ZuDQZnppB+CTO7wB3rILF5OgPUMa
WAfvvOEZ2mO8jxtwjyTLiWcfGHCHU2XXgrjaE/7fOpnFI5IG7T4DpiozWpc4C9OM
EjZgWwQG0koTnJYPp3KCoR5ZiO1/UrVcidwPPmiliQTzI47jJI8U5GcB5Gnt0+I+
4uiNtor1iQMO1W+yi/KpmUIWJsYXHh3zCrdIrUAo3t3/v46mziV/6iuL6XikM9D0
Skg84DR9+rXeZHGvU6AZjXUe/qG9w+8eZFPQutKbPDBgTnwN4obkSibGbg2nh7jd
eAhvGTMLhxhi+XEc+hy1/W5efzH4p74eczvn9wYtR8NWbndFEZaTl4qcFve3mBgN
KMVqh8t11SN1za+wXnPaU7OiIew6obDLA1HY5xu6sKAKh6kpXVNgeHENfztx7rZX
Dlq4ruBvc+Qt6iJvh7On1dO+EJKFzrT4abn3R+P6y4+v04SX5o/byX2zdtrLskLw
cEVeEC7dIDab3uY1hWWV1JPiWh26DDQ9kQVtlEAyGPd3wTk+xExwitDd3wIrQKcb
I8sRSLvQ6RmV07vZL0q1H8FKjhEtx84o96IL7IdkO1LqjBuqogsLAVaLsKDJD/G2
R5ru5lTxvqBACzzIdVpvrz4N+ShtUxZAWVcBHp6vQ2lyHGuVSfgad7D9+lniTCw1
ZkGRbgXdd7wuOfUBFmgTFoHsCT7CiaNFC8AOiBbenQAsLrUhknvqDGhqC3mg28w/
NSICL/Uhk0Z2QL9JwmepDFZFkMpLIZXXVmfjzfF7odQ0YJEIKPYr6yRlrqdI36Yo
Ou2LaBIvBB35POrl/vY3hfLohpjGlwr7+GW6kEnk+lF9O7A2tK2vER9LMaLgeEPZ
Kc2M0Jjipc5bCZzzIskrn8V/bcHFqAwjAD8NJCQa2Y0p1SXZ5wyMgyXI/DKfeazV
x2493x5uqAyz+L99DgEIjD4E5lU5xDxtMuPYewKd1MbXHSrsxAj7xaP0BwPz+TFS
32vb79es113frbalAmJN9dzDUipsHdElVuM8HOy6UJdrNBDAg6btU1zigNwVY6wv
Wj7V8cL5C+37KbgwykSlY6thaVgrI+mJTC7VHdJuv0ZYz58GDOXX7ZyDNHL7eUar
dXnzsE5tEOOPWrNRPASzhfoggM9Sg+kaq0a/16ZABVl4ty+Whq8EfHmkjda6fyRX
jvvj/1o/bJGoTWCt5sDEtBS5sVslEtqVKuo9EbjZ59BpWDabbzB4t4SIbViFrdK4
jwuz8/uXJL7BnsPl5M1vdMfWb167TD1hmBo8YRf3LYGzDGSW1+Liwh2g5WQxL5gg
bjGub9AKuc1u2u1mx1j16+k2QRU/AQkIsBsLQVjb04c/u1oJhC6b94/eOqolqrSc
DIYOFYBcii/1+fqyF2PV8BT+QYZtcynP051cJgBpXT524xN9yNCzqOzGpt9ETYpc
egIBOMcLRX9A/mHN6+QcgRZQYYFkonXcpgIbBJev4uUTUvScq2Z8tlciMH+HUThv
sdhDtOr/xdqtnDHlNe4uXf1NKOhEoEbstd74ESVcmNwFeHuFHe50uSH16cvyGA0s
oEz0CfHIVca0jaxsmstlZwjuXCD75JtwhhbvBFusoR6VkSWm07GnlLwiGNj7aY8g
W5m1wdFK1pz7rHOKFLQruWl4WpJV9GpipAsM62b+IRPrej24uiItfFSapD9dJ3jD
mfBjGRtzrxEn98b0PHNKJPMrtweTXB3+vXRozZF6TN6Z2awu1AV+Sf5ZRiwT7W5i
8e2HhQjHozWVvYl216bYbCp6KWV8qa2XbwSIWYDhm3aGI4KZffbAK0cvsV3o2S9f
i+xaNny0QwUe3dcNibIFel7VyRO7A3YauKAeZB40yvKmX1ttd19d+ZcMfCGlFbO/
Dac6zj52ZKkow1FQyRCyXmytnVbiku45ZN15f2D3Kwbj+zqodcK9gM5Bne2q3+PK
u2k8Yn5OWO7Mq/MopKUqGEwFXIGfsc6la/CPkQMh9qoU9LSzwLXt/ip6PkwXAQQQ
bfQY/0T9zotyohMr+wdZYG9Pp3y3IAISIArjrxJwqBAEOuTfxeNh/CXT0vELMh4B
bLELP9A4HUJTlIq6t9oU/mlgOJeJ+7Vj4R0SUZborQ5kEm2UuHX9lt/8KVnudmnI
L+99xSogZsTjgNMCIIbHXExWpjuq79QB9DdhEQZoTtFVubhM5I79XRmxn61O2u1d
p6vpJSXquZUkNMk6WUrBiWms8eWiglK5/7YUYvmNKA2AMsVK40kdaG4JrNC/p6Dm
byqrC2l/eHkRqKgN6JgM6QK62H59g6O71dRe3QdFY+N5Gde6iOV6MzKT/tJjupJz
gLh6u5QP1oNNbRWoTa9cYuod94E8sjzJYk0Y15r8VIxr9iM7KADRBU9L68x9NcI3
Lzq0TwzH3zmomd10iQatbotZ8VHHfiEx8aJPbkhbl9WnmDXRqIz8RlK0sczGWzeA
M2TqZDL4Ds2sCDz6+ClkgQFb4vLvBQ3llI78E2UER+U8dg9FnyTAvKcQNWT//0xa
mBXk1MsM83dtJ3vS1GF4DRNgjk2zlnilQ4XD1N+4xvTnKqVBW0+x63HrXyGjG8ZI
VT++9bzELPUp5IpO9jaaf5m75fGzWsi+XVSSQOr7Rgme2UsX/uTaH+wff6c34/Gi
hq06+0OW3aLJ+rLxOTUMjSahBTCKp5Ij+5S6djsSt7p3pQQ66zoU1DwIW6eRo6La
fp5ri73NuRcCXj4Q5bhoFZZWD5OOrkv2fjI9Nj9qfWdzhWRpDrNmKnCVExXPVKIH
zQRx3H0DIl83hVrV/TL/7lNrX2uHWjDV5Ks+ycNwYIYZDpwdtbk9zVp4wz64KOCs
PnsiWrSn8VPHrAH26EBpwA7AmxUW5vxQTXs21uo///sQcSPfqs8Dl1r8HSRrJ0jp
9/w9jQkV9GKS59ajhCI6Pt3G9FqxmsClGk9VoCnioDwO6CR14arRCsE3r8JeGJwK
d6CyftMaDCTIYfm40XZ1O1Q68zejMws0PSyCbr6AGzSmuTQqr42jSN1hIaZAoOeK
2aQ6Tx0meGjXqVnjy/gOOzjA0/V65bycN1yaR3XsXElaOMgc4fXsZ8brIMfV6UTS
ti9Lg/3+pQb0P83+jpOY/4t1/eDw3s8S3LSsMpgsp9EvUqun/46yqo2egS2sBgZU
5XLalw31otx9LD4Wkxp/nGXLZhEIH9+E12YkNRXjsECXxViWApkJWVVYa/y8AVJL
hrBnjWyzRpoGdt/T7785YUJ+Hh0+YlhbruBkDGyrB6crND8SgXk0H1mDAvf+oLcn
x9lUVXRFeEO5RSqJCJqaa+uhzPbgkbLDIHoBaNU8isgyMUtmYd2wdc/BRVY8GM4t
ePGbS+dH/DXSbLtGbliKH3UKTB0z0J+pil4ecHg5Vl4stoI/KPiVFNPnPRDcfXFb
h0U6RUnwRmaxhNJlrle06cKl2RuzxSsI44fpLYU9QaTmv1+Baf5/W4QyjdiDqEQW
CWoHE67blw8OKrGoSaPqVzLoGsNE721JXh95QshmXmG6geSnJfjOcnLQXbiRegzC
nu+PRHzFEiDjF5zLM3/tTXjpnlWOTTBTAnw7Hfi7oZ/0nPOAjry8V2dVi5lbXpMy
gBhXraBGsSAQIQbJN7TRbf3njdJSkpaHFGEEv6TDVCNW9laP4/X6SrOi6Nryoisb
3bstsWjKm2lRFS5yV3cditJLyjiyrllye5ymnOI57K6/P9442fytloB0h069llEs
/0GAkvb0OxsJP+xjHPSGXzKpaoqvIj8ZzI+HIgbxQcyR+L+MBfImY8p2ZjpDwrGX
0apAZuymCR+mbcuaI0Vpg5o+oT41Zmx5NL1hrrX7UZJQTLIj+l5kjqXvHsDxfVUw
U7+2vbuZ43zGwK93nQmYTj1aGnOy6khpG8LlYf16W62TS1P3g7wqgCPZdFcnk4sX
AUpsND6sd+7FisdtBPpkDzto/lzs15Jo5EmZXcyaEiiem0JZgy/h+xkXILCq+awC
+RadQ68L7oZe6C3lAX9TEQRDQ27N47wt00FAjCgifbIDMJmlswJuCmXHw1iQIDmO
/MVeC1VT0iRYb7TcPbcWMC0GjBpAWOPYZwnsxewxfs+TDeIZpvkY1jrQQjlUqnSe
JZF2aRyXsUCH/Mm3zdlnqT2rk1S4ytfFbxRpXHYN2MSv6qlU6LqOxauwCtzpZLqD
mGk1Lcps4yN44s1YX9bwwo0hzpltUUq2KeixmAqHcn1Wy+o/7Fw9vcrw6tmeCggi
K8fapf+jBwK1DOWZ9EFhE47Qb0A0wSD2ccQvbpQv4ogYJfxWoG9Rl+Vsr53D0+u5
fGSFfYBBGD6CfJ6UbA6nShMo9pB+hucqoal+XRc1TNIkUv3pO6NeO0xGcy6g5PCr
s58RoW7b7TMsUdfsEvRieT0I2+MdLIpcfCTXUfd79u4EC1cZh5JvsCY34B+/EjTh
uUnmzUZmUiThfo/OWWzU9438E3lpYWS/N34JmvtlNWjcJWsfQMNMCti1dNJGVUAm
vuihZam1rKQIJha08pcXsDVmHCFIt6AzsG2azk3XE1HiiXOdMTdGc/J8lWId2gay
dLf7DxeGk9k/N2Gwmd5kpWd2FgrgSAlAcZ6JjEVE8l39MvorQKEggDA+CgukRb5l
tV/JnV7v2NB10aqocWM8ZQTV8hyM6D+KvASkVTylHQIQLLTuZOHUmq4vq4P8jNHb
gQ3VNig7tbDlBhFfREnkrmStfShI4/Ej/dSNCfug8+0uuoAUNFNExE0rF2vsm7LT
O9YgZR9/WgtFXkIc3l9pOrr3uo84jas4Y4VRht/I1neJeGsmpQ5rVLjqgFckoBCc
0v9Czqv5pJRet0q1P+JRhwvomCvOmWtG915vG1KOlFlW+VoNS2rhNg01iQUYRUFH
XxEu6yMTHxp4ViNjDeYMK7opQe/Yn8ltUgns2FXE7vedO1YC38jOpo/blqRt5/V5
1H1/VaQ7idHdJCvzyyiW3B9FuqOmXnjFISL6BxGMuYtxkIsBYd1fojRDhSd9etY8
85yCXBAd0+a3mBUevTwZtbZcT0A5gDVSFQM4ymaf+1e5JHXtKy0Q/EQdqyCucc24
H6+tR2FAjkgb1U+BGmTWh5ZlRG2UfdSuXo7QzCYnd1QZCGi/5fPArCvNt3qH/gqD
inSsjiCPwbac6lW96BuVWllvBouTex8nZ3WLwyPtw3pTDxlrzNblgZbe8dOf/rJj
n2wqN2SVqHelE7rYF5h2NvGYeiRvHuzYMHgCNrPoehrYp2XAM6spEtEZbCV793GM
fLv2S0iB3NZyzY5mD5j010/04HBtTUAqyZE5K9I/Dktj2ZdUytWtbnQvd8DzR2aP
+Dqs3yxi4TnvcxE3hdvNPKCOktqigezpJ8SU7xNGuVHjxoPsLA85M/dcbabe2ida
+SbCPBll4dhhFpR/tEnnV6dMhMnO4LRVEdtNAWCa6WXQkYekEGy1v2GfoBrJ+wZx
b8PtPmACilFj9qZCItFIONX+2ssL+/Srp2143+5AR9Wpi9mM5mr6x4rLAdsF0PEk
ztA/e9uDymyDrFyZnNg8dJEJ+UQoV1r57P4vuH9KhMEqzaJ7bpU9Rm3gkl7wk64i
wOLX8Qxortf9G4+CQrqC53VaAe5juF8MBwuoBrT9ivVRWME+SFI6TE0P6S68l6uJ
aQblX1n4s06uNXWEkhSeFILNkA73kNmWeHeU2/GrG//Dn4hr6x21vKN1arCbGGB7
gJZCQpBfnDvLNNkz6+LH6i3A8QBItV0n3gXuo5XvoQLllqce2TKu/kk5RQykn7d+
3Lolcde76O3zpJ7AhzyZUAvBJ7HeXkRgJc/ffUEk7QEQQsJuorrb1flqZPpmStvB
ztoalEkbyNZbyKfePQ/GRXn53fVC3zonIf9NfLP8G7ERdo3ixIgKImDh+G5fGdnS
U1IJIYPgIPRO4+sApZR5WJgvRAan6ljN28H/I8Jz0xi0nPEFnqQLx0JVt6Buul7m
AgHp1iu7vUbtNDHGGw0cv9enCe4JLDbwk7UITokknZjbHIUqmrQYVD/MQELJphfK
4gTzElVh58MBGjQNoBsK6YAFAOG1oqof4GuNiCS/sAYfWGl0nD1vbZd4SmH9D6Vb
PvObGPSMmM+e6gXbMB99Yb0Fc718xZ/MGer+ZY+u9/hnjBo6j1eRb3eBWUd0dPu8
wfM9aE2LmxTw3RAV1ii4CZIwCE3S6+mTwaonTbd+6zAu5NDngNuw2cBVKFGt+C+D
gESz6rIA/bkWGr2fHKsg4ZfQEXuDkfMPM1nYi1RusGG2p11EJtMN7Obk54YToxN1
5dkx6LbmEGmpGyRWATtQtqAHgjlAGrGn6Ep0CU7QqxkXM7zhul9eo3ZwxbSFwQNu
US3ICc/SXTeolvcXcpQ1opW4NMrJMq70+uBsdhmVBn34I7IxrYsHtbFKnIsAxXtv
wPL+zz3jjLbZb5eNngvBXTitwUP/hJkoEzFkQO/mhK8gcz2jkZhdv0wWmcCI6TP3
WALAOYld3CZTf+1jBmc2pCd7wlGwV3vgwip66Rr+22X59ywjEt1Y/6C6/leC61t6
aof0Uxy9OWPouPVz8UpHU8Z2q+Y2yBLQCl3o1/pq3hcqfMOPKUKslMKquqDWgsJr
kHV7fRuXttxMNEoI+PHrzJoA/1BQLn/WRDoqJRrQpxJhVKDfCNMiUJQ6gmcAifhS
66xhrVo5iIinGJ+EkBJP1t3Hft4olooa7AozVPVm3GaV9BNMrJFyP/UXeW1iNrTY
NyOHU6ZCG8gySpwIzzF16WHw1en5AaIgFyaP6GSMZ9L5dKVw/K1KIVdF7OHidmRE
viwkPo+SZqM4csaSsSw3cBFOTisbUmmBMVHPEJnK4RIcjlWD9CjeqavqYuPxOyBt
hkzFHagFUzu7FMhGCUaZA+/9ZS2n/8bRyS3OtQV1TNXs7R9EeCcKG2uXasgEucFw
UYP60bYf7cd0V6n/wXh97bIUQVvNgM+dF5vzPx79PCKoroAcUX4ByyAbQiUWGLQv
pNgPH6jO0/oiSXGjaF3FBJ9Os5Q9Nw23aBWBatLmDsCboQ5AEy5E/3724/s8Gxi2
5J12pIYfVmHzrjYR0GhaNgmKKIcclyljh9Oi0IhuwQYcs3Map9NKayCezuhCZOXw
xA2nxuVyA9l35IxcokOAD0n7sYg8s0FWFE8WkjyJEPGXpdTXvJF/VtWNJnIY1SSM
lCRjdCp8kW1Yl7il0DvQv/+GMQQSOBP1kNGRXyJq2v/wayDVk1QIA1GALMeS8L0N
f3W0nl9UcWz2lWDFAeMVwZhtPw/Cj84EOyNf3gcd4dks9zjXb98nBz6Vms2sOwd0
3TE4qsaixef4k0HlfDN4MwmCV4edAJRINxxi2amo2RBhCBcvk0ttjL1AF67yylGu
QglDGLrTKzmscMlB/YAxE2KsCzSwKuoU2fs7kKP/69m7uOmQ5ZFNfcpzSNCQurw5
4gegltfiGTmxnQ5WH/r7+knPgWijIBP+ghx+1aawClTZ/E5tmIo/zofK3uUjokP4
ZLSaANyQoP74wmzv7lgNu0GJyaAjkJcQKZBE6dywM52qEk/q134L3Q5RJXesOPcA
kBTHZ21mDl47ffNsQdCXYnb/5Vjs4YQW12Vl8JJSb6Q3GW+CacvNWfc1p81tC47f
k10ihi/CU3xkOEUsRNwatRGfZuaUPcwukl5xfe7up9yLuC7i4gBgj38FtX5mFD3r
BmxY+nsejVR+P7WdvZCRdLwcm+tvRfK0tfRJeDUwCc94KY/xOTVNGacLGAXqWOqY
CpQXg1WIeQH5lNQnA0BiVncPb4Nj51IwV/gmAjP1dSvzVQU/kiNiOj2dPeCF0W07
rMInVSlD8YPHe3f2bo/HHzGGKs6P0N4qSS15GRfIkVXHkab+A+Caw7mB1GuhstwH
YmrMdPwPk+ZZbLXBaUs6CIJ2MkuwfLOn0P6FKW7hEXLAV6bGBZ+J1y0wQswVhzXH
u4JgsHLuVEY9emEUXs9DZkzQRdYX7Vvl29P0NAZzgsecOXDUNEvPgPEwfczR1oxz
wnJlDpm2Yxb0GrpQ7myjmkMsv+KkfELjwNw97iEp0SyIROmfyIR9WNaKrJ+2JNg+
G7pnLfsMasb9coewalMBVt54tBQRmkOHD3VRvN2Cfj5fUK2oauSjyZi/3GgLYZaW
LhuGpDdwzPYNpVTMb0DfzS8+hgvA38ufRYvof/P2zWgQqbwZuGVu+Eo+KGAL8bVL
SEih6xxMt7vv7SdfKzcDcRU8polBBYMjmrX05b61rjM7oKyKz1Ms69FDnr1kJuOL
WFZh6XqIOAG9h+Yum8MbU6N/1R6BUCZMOAfenyD0CivwZqiVRPMYJkONZou2PLj2
yugWiVPLv2Cbcag04a9j3HOvNi6mhF1xtfXK+oxZ+j5hpSDHkyxtemNgDkYACTE0
EXxONohLQL6w1t3V6vBtpaAe4Vv4oJTFhDu6/fzZNmYkcfGLQrAUM7QqmW5KtaAg
SC4A5l9oPCRR/jEsoaRqAy++TkLUF7Hfb7cqSdSLRC3IEx9CixoKgzwvIOdm9lHP
lawgFDGLgtz6pieannzkxae6qCyoQhqtbgyZc67JeqruGSVhUJt+Fl8mSP4YOZVY
XGtrVBvTIwS4tWtbFqTMO5TnhDdNstJWyigkVR8mZwKvtp/BqHvWz/pJvOR9Ef8W
TfuwLPHNhzK9OlgNAK9rEqTYm6djR06USZI77LShXjeLRdKBcGJTzuKfU7k+K+2Q
wMhaWXUY2jKrIIej0k58rsq92RDDv68T/vGi8Y/zfoTavIO6mxU3LWkwh1J/IVEn
GppiXbFycveGGvg7u+LNql7HOklU7+n+TZlumt0jAD2/miMWWmSzC8BpD1CcKwC8
uMh8/A54ejfU12oGe2ADU7OyycVo3xT83LNOLhrrBuccvxNj22qVIbyd/Sb151uE
FgPLebhGielBQPTcHWzRCgvJV8IbJltXulDPJMSNNJQqUcRoryiYxHJb+B/LdTLP
Q0/V5oGgoLQFFYpySYh6dy2je4C2QC4E4DdfyXsqK1NfRULC1afjtUPDycKR+mkA
D8Fy5m51WcOCqXqmGv1UHSQ1kdfiYiZQ4nzF58m5qvR5YS2sDgVtSesEypokg1ZA
hLTuEpswYOhQKEDAOlfmetLngVih5ZgRg4b/SW6za/OpXjzPWIy+kbBogRBGjUQu
O7bogH7BuxC9X+gBN5pqP9j5amMvPuB2yoPGiOj+rT4wEH1oMSMVhsAuWWMP0tUN
za49JOUwoFkdHwkl3mGS7xtzBBHSQ96hyDXuCnBKXf931YmcJReTjqxANHNq6f1K
+NFfeYPcA9kKxUMRXSyOYHPBYz+C9RTB2+gErvghM3937MNXc4tLHxO73m5EvClj
EMMwuyZOjL84r2rBkqDFH4wzm+geEyFGfh1+hZQhyOZx96T9mPXA1Az4JjXuP+28
PvhT+o86BzyQGPMa+uiUJkPaJJLHhfts13vY9xf5JayWknGTohcp3q/Hb6UZwdhX
F5gXlosobhiN3l3WjSmP9G9Sp5jZBuoeNvbgpm3/fMGUanBGmD6+RQWLpsBk0uqO
E4P3SE8iYdK9Fj8HbkLwDzWx+yg8LhWgPVi391WJaNub3o/NkiqmmxUlE/1a6uPR
zwLiEP1fpa4y5uUNY/CMsVj8QtbBiK35XC/er1arVVEAVzQfu7WgIjzkeAodK1a/
vJSyEJMS+2tA9Bvbt0dUsrg0qAFARdOMYcpd/N1EgDUp3K6UvxP9omZKBesXKzLb
l3F4cKSXUUy4MDMy14W3lVRxOd9UuxrhhR1Ihu+m0yNMGEGO1+pHIfza5msRACum
Gr5ICG9ARXwe2DaZyTvXH4H2ovh4mxFQxELkZffQ+iCu27+uiuG0/fssw68WmZ3P
mxkjYMu4GujW2V8PuOQUTxZmw0ZhZpkuZWTL4AIE5yrXjmFifPwlYwzfY+TvlCGV
qHgLYdhZhEKwX0QOJixRsv8t6tOdDn1zN3pyflg+sEN9zhkjUwL+gSIddYkMC+AA
s+z1bLtyUc9JJmFTlyg2tk6qldw+e9XwNbjEYBdHE0us5zjxqto+3p2Vpj5WGEQe
ASsE3BxyUk3vhe25MV0EO9ZeFnZ2PzMEKeh4TVynTRPaMprMjqIccwD+xOOjF7KZ
suduwVqBz0cmXiLtfbXK9VtwaJy4iNiPDN084Lm0awo4idiA2EjraxpSXOoymncq
dyDPem70SvTFjig/mGMjCqwsl51gwZ21bs9TCi1oPXXO6VYxATbXGybQ/x+JB3pf
50N06WrfAjK2a562Mhm2UgV7cMFklYN3JU8tYgWLEtph6qir24wP6RkGcK2rFyWX
jRgWCNhfwUQ5SHnZtNoTkoRj3v+zRu36gaDxXCPgwDWOCnMZ4P8IiffRD7N91NEJ
4aifg/9wlHfnMe08EaZHYQi8kcZozzTwufPyIY3b9NiXVtpf/cdEgaCidf+4McYK
fPJurIMR9SgojEuXv5eO10KNUmefX77RSqTya8new/0VVoz8Ec4njcmAT6f3VTOr
qSPluiKs7VMytEKzWKHrKmz0suVu++8N/4FZSg9Jg46TR7zBVOuT8uVby7uVG6Au
QtKIOOdL3T/Y/LA56j/F9NzbNkPXsRkT08y5H7UAgR4PZ8A04QQlfZNRvO/051zG
oAvRoxXG/i3E6vRAwJbR/8E5OzACMFTku4ZV2674yUR2YnskurgiYXc6kS/udKey
mJdorjIg98VKW3ZqXYq326vRo731noRB6Y9KYbUHnpv42EZ/WTFGCpDX8u5YXkGx
K+/KHy/8tWXFImv5jEmkDYgzH8dlpniqQKzM8WnSBCKpL+hKXbhwKaZ2HEHalsUK
xVlT3H9kHdyNXPCKuhNPqbvnTneWYWsjoI6y9iEfdFENlg1PC+qbO0WHYM18n9+d
i4I+jJJiy9h2qAAjmYiy8m430Ri79sXokzVXl8EBCeOw4vQpFBF3Hd8MxpGW4ADF
9qZT7u5QRyh7B00XtujDtZacn/+UVCv9zJ5oLl2PR2EPcbcGZDKyzKMsceJ4f8Bx
dasxKlTvi9zbvoIaBkpm6ISG61hfYuHfXX6CtEVH00y6rHqTlj2Ud7EpE8Q3meKT
lWw6j6LHPecwPf4oNiKZl0UbX4lvZHSKvVDeluzEf6BksgySnJTklhU0rQT8ntzo
SQUA+HLmNSfS9So4ZnK5jqTLMtu5uUTAcfbAd1E39jOIzC2nbSKwpqdazDO7gRly
DTVOUStJnJQlmJ/C0u4daYdADroIPTmXw+lYLkZuRrsNj8xD8bZefO8hIz8Vc9EH
EdvrZNgYc5gpYY06J5F0iR4MTByZqCXiFVOw/wqR1Kga3ulgqGdL+01vdANMUNpS
a61SY91pg24QyTEjdyWZETV6oK4Xh4L1pAKlBj2tK1F8OrsgXPD5q3y6id/NYwIB
rQ3tlYKj6FIC8fY1dxL5Stx3YOxa/IX2apaQSkYM2s4nmZ4RnVNNnOBGiV4JJGbg
cjeO5uL7OJderGiuw5aXzhu88l6r/wDXnWeaZLOTwcpLuXxIdCNCDBrEkls0BHJq
wkt7CCJlAZX4+aC720Gux5zxRehgF6etN4/+HmksJKG+jmwOOq9Ei8VcORGyaIKu
aDILdMwL222TwtWX/bQ15Lt3uJVIqtNMnuG7donMHrOfuitDpEbqHhGec3BIFn6p
IYUj2JGPfw2lYJMab+74V98kZciZGWbRGbGl7WNemjevZamyM5jKB9lYnDx4hGOh
G/NMgyEmZkbtC/fQMfTHJq/KlIe8fPnvSbSgDC2GjeHtdghawmZH5ZeXPJl9PTJG
dyOJJTlR2w2fSmGPbCq6Zf6T8IDk6VGUDfatr9kHUVhGIIMtdAigsjW460Pny6bP
fwO5xrzbrbldFSnSCvhOm/ivcS9nXhl6gzdKoUweNkpFX0knO1tcR/0X/tUslvL2
P7ehIGjRsXB8Yp6yziweMn8E1fSHDFCnnmsLyHxjlycw7M0f30TwukpLNMQvConx
m1EAQEXp04fnC4B6cPlaRg6RJkaYF9k6VCHmlikb2/oIj/1oD0VbLw/NWwYjnqIP
6s1HDHKK/qMDeITuIhizS5Hmz22yxS3HJmqkH5tiWX00HyzxuMn9bqFQpSvdEvxk
iIVOJbYgqdUe9QNxd51Q80RUxtfLWbhoaFsV0L9+av3N+j46EF3ixbCzzRArg+PA
TWYyoIhXXtI/QNt/IsZ1SDXU6SNgeXfhD9EON0ZMKTDlDyWp3dZIcqJFqBI030rN
gOGbrpS+hTncQr/1eRiYej8VaJn53isJzZLrHn5TXCtdTDDWzf8jd4NYTJK/+Utx
npiaT92pjo9oGsXjOh2zZJIJSuZd9RvXYVYWVI4n0+KXTpbHcfeuSR/wuTcyR+Oq
tott2khrvNQ9ak1YTAI3bU82152VPWntAnX8yONFCNJXYpFH1WOHL/C39G0h+kkS
KOZ0/2DjMw+rswWH5psTWnw/UA3m0fdSoQ6BrWO812z5QIZQ5tmt9JWKvSjZwePI
3fQ9FCgce9p1TtKUP2AIwPl4r8hw7Y9nhEGwTpgwIBXwpUWdBPV7M0gHkXHBKyMk
j4dhFLqqhAt3CWDVm1sLJUPAGVXlLhwhsNsMIeE2u/X2PfF6wnFFRMWCvr7LmtgK
KuhvvD5rnL7bQ5To6/fW8kVWHkgfTt4gGKNzX7avsbBv7PfbquFJJFv9YYOXNzb8
GyJmj+OtxuKRNrmievs4a/mMCHJVJNpok2EMSH7Of+lks1iRlBTOcP4luEhQ+QwX
NB+SeFXuQUBCXT7/p2vxmgwuvbPBYcih99psmaf4LTmMRJJVQJ5fGMxSaQ6nstU3
UmJoLDHTgxvZG8HFSQ0n//2LW2vV2C62mD4iGOwl4kpyFfZ29kO/94Ql3OWcz9ir
k1LVpFx0CW3tbEW9j6Lkpm1Xfx+z6ICknTN2QzB0zw70iPf1dsx6k2ZSwxviu84C
PLjziZIdYASEf3KXb2YxLe67Uylx4DkQaAq9IEO5XkZSJaDdTkNd/2U3kyd0Anmo
qkNQDI/0P0JUZID8gLBjhidzuFAcpYs10huNVhnv2+tzwFNPkfXbpyCwVXXpoTnu
r9EeMnNxqVLZ+rWsXbHYlVaHWBCqQi8S5XPg2wFn65VUjFq3MkanSWhMaRUWDzvC
2qTjLUYJ8P1rIpK9b+cOieC3/2D6//6c0+E1VgF1vHQDSVsibNf0Wtzp04Qq4bu3
RQKdUeFCcZfMWoiS1F5PtrjptDA9v2rUQ9xVVy9LksAcUo7du5/6mET5lqtV1HHN
N1Ya8DajhXMLR36qwn/WGjAdKX5gAAwnai3YHrYYRfdjW3NK2LkJzezVFt+vlmKH
ILHGvhm3maXY7vkIfk1FkDd6sotgFdceeSSwJSrtbpwY/1YdKYkYSzKYwu6v8oLP
aF3RtRSr1QuPPP6XUvLw0QAMLQwdist3jAyjld2uVPJw7kkAml/nupNEXe6kXPsG
NCzYUG2+dTlgLyLL3rD6cmcoX1cbJJ1zJpOy/9+kNhBPgzK77YhzqPrIRTrV8wx+
1vtOa3Q/9goex0uVrZCAMn+fWgbhimXVBGvx3O2mHGpCEcV7dFDlpzaRPuc0cZvS
F6c1h1qZQd8nKPrPGsudGa8W4jlH0vfODuKixg09MqtBTsQwakfscApesOZS5Y/k
/5bLTS8FPmQc3kZVXFrJnmyjMsfbkDJVD0dGJsJb+VJUTTtOuWwvia05ooQd5FAz
K18oxnqVk87jtrUsosDQJfDcV5DVSrM/D9cvw6j7QkvAcu5FsoQKpg7luAz7Axb0
vd+gJqaSdlZTSk8pl5itssed9Vmj9gQmAFXQgNIuhhVcm80J7VFINNaCEBDf48Se
rWxtFHjwCkwan094hXcXE8QD2dkLHb4uRmUq6dY0m2ckIvvnu6PtGCsAdMtSSjCY
Ojnhj1ALQylGJeoMNDKbPAmDyduCYMZwMpZnlAIFRVi1FzJPU42num5tZtQg8ytk
JawbhR5TTTje+n5rju8aKQwvOUBmxqpJ/zo4SRbU5vDPvvSwaEYY2MaxskZFOkEW
cAOArs3hLk6JtF2jkp6uSgFjY0rT/3foybzfrUlj8GJNKYpwwvi7iZ31Pju0LPqh
Qet9cGZaSyz62GP9Y5XnyRUCr45ojgBvINyCzLxE+F5UGDWOrdaJ5twiLVdz0Yss
Ce68m5j7QGKA8Yd+lNJ6hyhXFX2qKELoCPl6fEEj91k8xKFhLXJMcf9+a/qVm0pO
9Y5kCPPuOeJ6MPJI8puxzTeUrDSamESwqkYSVohpFCITdLMdCWHnnZc/mlH8DyBM
W6a64Ror0kZpqxpnzIdDr+hEg3bC5l4fGAMVjBRkRVXLfYOyDUEJnBp9zdwu2JhH
T75LJy8HzCSBGCqaD8dclJnl11TnIlaP1e73x7SIqwwSPjxWFw/SmboigQi0kmCp
lJL5KixosMjteOGvY9yNEseiL8iBxGuYwQJbJ9+UY7e++t3OBFMapNycLlR2Y2zH
1XHZXYnbB4AwNnEOpl6keUreidTT3QnYcKdabs1TQ+V70d7qWUDSIOAjjs3MyZab
7RbgLEfRlbfzS+GnRPPdoPM9UHmkzzTJ5kf2c4p+7Uouuuc3uLqRRZ0x/xCnXIyo
O15t4q0SlcqE4VsUlPIg7TVtl4fEaiouM7OY9Uw07FfeuiJLypV7wIvptLP3gjCb
xNYvU0/hx77Pch2ua+g/4MV3NISFuqYQuMxSE5zTVkZmxhn5YO9zf3cEY7lR6hxP
J01XKbzstfRF5z6q3HmK9VwTQOiBelYBEjJRVD7nfwexfx4zMD3PE6fhYm8Z4LSq
5IMtT5rOPfJpyQUEfKdgilmgDFKRYCoUFiUx5OwCyX69Ry08StwjaWFosSGuuOlV
wnrKezK+EoT7CVxfDLp+6G53cz9sONz4wYDdamq8c9rzZyAuCAH+dA6pE/sQ2Zaz
OuELgL0bq6Rk18R0uwA6U9jXdjQX3JbCTB5e5UrHbJN0iSkTFZNIPIQTPd/IfU5R
akoawgRkcH8w+QDHyGfGs4IXYOsDxcm28riN+n5xSpxohJxO+R+yIDfLIvW0beaK
ksuQ8EiwWb+vUNDGlVnfE8CsAoW5PKy9wNqre80/MbVzWRn/sCiXJf/g++2atm40
bnEtznChCgZ50jvmxAyXeABZsT96mvnDbW398GwhMWe8AmQZJH3Y3ISXtyZf+2GC
Nzs+gvpm0hLvNVRq+p2hSN+iK4s6JJV53iZGBnN+Divb8CALkKmC0FK6FP6JiDlx
Y8dQnS9FHClAZcAL1+hzlwUCthlpin+rDc77jBo+/We/fpg0OHUxAiFfdld1Ea2p
bWdtdDxj4fEpZxzOeO+A6gao35t+1Q6GVMP8HJyAhnrWt5y347zHlCSrSvLUb2c3
sD88dGAcq97IwRGS9yZiAu3n1lMghHQoSIhSR/DBbK4vQYtVOUO7gPjznMcKfgNS
TUU9Oo/vFsIInO+IbJIn3y9myfETYOhAJ62iDjoHq79OOtMVEVKDIdPydhtpreeJ
bpLTaLp/sMylGOoc8VySs4zgQa/6sGGW1nD4CtYksxjjxNEopBeuJXlItNXwMQ0Z
jjwxK7sGq4d4fvSl09PGH0VQ0SVqr+d6VxRbZNRpYbUrDtDQgVQEAHsu+9uQf96i
5DBp/iHyNMfp7X2izRtrrEln0Rm/WCvvgCYr2ctdnjCQ9v7xlzCSTX68U7kndEQr
jZJnxGOX9jdYmVbQ5neCb8+PNSSE68DizjSJ6pxSjS88SQdgyImQan9ph5dwMPbT
/d7AlaRQLmgLTw+ynh694VRcys3Lv3kU90TisLVTAXXWzj6O9Krtsx9k6dT4UQIh
0RvFMqDK6ZDgvJ/Z5dRuy8RnBCBCABaT9pUayX3qRMIeEm85C7NItC6VeN7vHStw
GBDIV2/Ufe1iC6bznBFQVkR/jmOHwIb0EKVDZbGQn63bxnvS3LMoEd+zFFyyzCae
9QHW4F7SdNdxTKjbQhwzSseqtn/A3bbcQUF0/k/1v725gvYEvj1uLD/YIXeBZY9k
+s8XVitFllPbB3+L/leuGQ/c4NefmwlfwCbhtnrWMn426MSUSSFvhO3mHFACYlyX
7NrysKc5w2paPngFnkpFB+wGEQomK/DtvKEt256dVe2TJ/XrjVG4wUPW2xheOn73
mOqGT6t3DTv1t05252sV3+I5Xh9w2ZPRECnH/FAhiwudZfPnuQthQ2sCymwI1v3q
O94GgGCVXf4KcfSOZx4JcM3BHY35s/D4JAJ4xF4YS59Ea+sAqLj92UyrqFVJC3iY
Lmj28kvfNPI3oAU/juDJLJQBA3T3UlcTnVGVPMN6afdEwlrN8cG8RCfRBkaH3PuJ
gIl1QinafwCxRlXpXl1SMMR3ehu0o2XC1awDALNVyhWp6tJSBjZPXNwuT+zQSmAk
OA1VAVswRFvefuQRPjLKmb90CcotdPux8uYtM63Fg+KZLO2Fd4ePLOm9MC1PAFhC
nMJzVqKDe2k46k0PIOxvV6hQ4scQmOs8EmhgmgMqvmyVgYmNSJA1rn8NPATFx8Zs
wOOnA5KHytareRY05u7/5fnUitN3fkzcHuIsmI8j9WcerX3mzRxghkyFahrnznxH
DXMQXOmoo37L99djdATCp4z+3ntdfVKIxG5LlkMSvry0/MDPU0WEwZ1VV7BZkk7X
iQIi5A3xxxkNfPQ0waG1VQ5lb/WFvSKmMHvJbM5ST1pa596pUdMGvhM0O0lr7d4Z
K/2QsZtjpGhxDMwHsQXWbtgOrOYx3eWUkmazKj/fR5mBVLXPk6DSEOZurqb145II
pA2w7sut5wA2VmYmWPZCxD/cDRMGPae2wuAR1+w8fy+M7HgW6PvsE1AGkzrWMINJ
yqqs/Qih8O0GyB0+1PnhlLorZFb+6eShFhIU3HuqQUIDqzgjZhGucKhqBLDq8eHt
xU946j7qxr5Y5sMS695cVNuqAFieOtqcJSb/P/RjC/Tym9oTjbSSevH+8ShbdGKs
zyiIVkpygWcCKgkG/0jk1NEmW6XXaLWRYFCYVHjtgpnzAb0CmzFZ/q5rbvhsQWOP
JKyhXHvuSV1kER63d1M8ThTqzlLRAGzpHaoj54F7UutPRwFZtFjxOTMp0gLu7cbG
DOUMyII6l0RXkXIUOBjNtQ+JMRZezs9AH4vh0SmCZhouBBMoqpT5brkgeFtCjf1V
K6J5yO2Oz1r43gXstdHK8Wh9HNgyc1imReIZ6WlCWnHFz0nAFigXBQ95WFwxsV04
DZaEyuLX9fxe4wNXllDnTdNDwayy5Q84DSsA5iYCrjNat2TL61lRo1wKg9q0/D/Z
eFvQZyFKc4r11E4XLlE6cjlvVM2tKbijidF/TqmurG76z+zPr61o4nbPGDXSY18I
hoFgXF9npXcTnA88sGWwbxkIrunUrgZMcF4anspj2FyfiK4guBYb+wQzbySdWIhG
Q0qnNyMRt1CgmvkwKF9MGXUxmOBa0imAC1v7OQkXHLag02ZPlqul3kKfcdo9Xn36
gTOCu7Fy/8Z+H6njUx470+VdiOyTgzO0dSy9LumLRJveZxN3UKx56LUsryS58RPR
keyB4DyLibTvgYRrKuy6O+GdnqE4Wx1erGOh7tgK7Vqh4a5em43PxoY9N2ftYhpB
7ShM+sMN6U5x0iR6gS4F+a4UTFmMJACVFARXlpSg/GcpeKfUfcfLTF8Lxht8yibb
LksLhP8uA1cdOhX4A28yeMQz55Bs4L8i0PPMPeiBuMYZXRe6CQcn8fFqJTKJCykS
IPQO+LRxMPFnweFj6H+W84qJZGqhNeCV7tdVoSZB42ronrZahhj8lF/6RjKbuXyv
p70Zh0odifbM6qOJM5hfKee44NaRTDLMpkMnKJFDBbwjGKuHvchrQPbismP7461y
AhoVfF7en9oxcH4UdVSXOzXWXvd10nfgGr4Pbm3lLuDV8WHFJ1zNPhQMMgmK6Upo
Y5+Bh7viEM9femNZIcYOLSHnc297OX15o6ukp1+wTwO8h8JBfEWRLmHO+54j99JA
e9f6+j12ccmt97rK065VkI6iaJT4trxKKrJeSI8RZEYEdnHAM6gfbiwBmFKEP5m5
o/WjMVC44trAa0U2ryBHdf8mzFyvzV275Aot+1iN9tyQTq4sZa2jWI3KvTY4rLml
lQY3yMvphi0CPjWGyCtrbJAMuyRyvdF2besL1kr0XpC0kbF5RdxZjOygcVW0O9JV
esPCR9/qUElpsy3ZSbeRAHTuucFqpZ4+GwNTc0lCDtoA3unbtOWoOPnZui6ML32V
5I7lpVkiIIWjaCxV/QJaI1jO2TBBg89XEq1t1yN0CG10lOVf7d2grHD7qkoFGkCt
FRc0NzhrunUl648A1zR1+BH1UE7BZ+jGs1H00rfzaLIISZ1HydYkPm8HcdqLi3PH
OlnWosFXgyllO0pUxbxgJU9V2Ec0NFqEMByy0eg8330xql6G7tK31t4dqZl/UJlb
WO+OlM+Qkx5+cN+p2XyykR8Zy4sOvyytE7bLr17+j8hLFvBYfn8bP2Y5IiH7dEIb
r3qeqPZuM3uvvJ/EGrAhT4Ss9qEN0myZF+J949vLd+UZticJELLjbl6JmsxZCU4p
/pA7wyO6nbFWNSotXrFDqJgadcLHuetiFeUI1atwStVbx1Z/CstoE9WOP5xPf6JB
tDCfoEuaALyzM9GuR5Veoz0FmaLUsJNxyMGkm7uDi5OQtGYvT7R02neuW60Se0pC
U9QpDGyg/1tYhkIRt22OB3lY11ZIjIR6+o2UXr67XViMwXBHxyMrXLnoXiPy2mVB
/t6e3vMAKlLrX0UJhCXa8cyMzs9SwkW4uszzjbzK12uZWpFKBH4gnBbo5nTyPZRP
0XMsH7qWye9Ikw09fzIO5EX4PP+6znBIornuPwgNU0TsWCb37wicbq207fbBOQ4m
4QyRNpkm8L9DAN2Gd4/MskI9ewyXiL8NJJdTp2tzv+1zqPkdsNYR5hq64oxiiBNi
uCXCt3kxYrnDxKxYVLYjBUCBb88mD5zeIIdIoCDPsx+FnTEW36JPPo88NSNJqzC8
cElN41J1pSZOGK71K3Zcp6pwZhSZfTWhtwfDBwvvtjpDUFgSlGACOAj1b3DUtXGY
a/vx0MD+rqFBKBickQQ7mQMkjT5cUdYzZDmt/L+C2uQqUynAy1yh8po+4ES+VtMH
9XZgA6Tg0KpcCkcy8Gsn68b+ab2NSW3+w1L1u/km3MtvIctO4vYJIwb/KAlJXDew
CtdYGO7VJL2R6GpJsUsZIOCCR6xNRE5lTSOAmMdSAEI9uOJHUw25HiYMa4DUqXA+
o3P/NnpLiX1RvKhpmGS8zpRXCQSdMI83p1RTeellSybnelJU1NhpTI+kAYBMBv4E
nGge6vDtnetnIUaZZQZyKlwp8r0EQ13sEc3MziX0KqLgEiWEfsvlCAXSzXh6YoW+
bi1kb5l3sePcUqv7tpMo4ss8M62FRbc4zSui03TytmCyfBzi2wYJVseSExx9eXKv
J47A0VTy8Gz5EORuOOEadwDOEmBXWU2p5C5z2IAk8dfx/jR5ct60SBTvRR80g/Xv
ffAQ+a+mYVnBxlDAi/s8F1F+HfAL3XFQwrgAcRBphZ89OfqYBR1tpA/yhhbK796E
oAhK7LXqyfbPDWN2Y3p1akEKYoC4crwoScrFH9qVVB8Aa3ExNUJxJA+yUup0jj3t
1DTQZo51ZxrhcjL8C0JhJCaOao2dQwUPDlPdHp/VYbVQEeuri0Iq6oAW0F05o3EJ
JVb0zD/QhbYKMycBOOw5iQrzTlCCJYG9Gk2hmb53XZmJoyrlIKcpTKYoEeHpvB/V
IQelSYh5h9wCO2Edvo66jWHP84mBZcjTLqz65HLIqvz3ni3qiHO4+Q4fxxAdwCaG
b6UVeFhMAOyr05gqq+AO6bylb3PzUPQ/XFhMP2bNHYSFekkN9RkGYeXUeQNqNA1k
86IKrzKgTo6RUFeWHUn2rNIPiEWJWYjsV1a3Ffv3+QE21VJOAkpqk0Oxjtw7d6Qa
TFwhvoIohy9z0D4qrnzSug21QMkIqYzyWgUDXQIHL9kfY2sgmmybXY+S1Jm/itSH
twM2muchHt5mmleMwpI13pPLw24xKnxcPFKclnWXOq+lNwgBZd03HqFSEfnq1yo2
QhxzVJKdsDicoHYq3k4xkfKxynyO23fibAF5DYBdqCd3d2i/ON87gwasMhuyXiU8
jlVvmjqg6v36mfZuuoevAAL3rtmXc+YDWymN6LDpJvPPd5IhXQcjqoNDFKe1n4aL
3znjUmWKZgzGnA2GohdxgS5QaGuA5iHvIfw7d8+9Mh64NAl5i/Db6q+dfJw4wLVy
AP5bQntSObBa2Feh5BTGAhmDFRcZGyRcG1A22qeJGA9OhL3S4UnO7ikY85hZYwIk
c4cEnKbsTi1pHmdiEPjb73NdPkNk4FDDpOz5VGKoNLO+ob5r55JWsRBVC196Ebh6
rsqspo4wJvMToe52OvAR2HKMvCGxVuO1VHmuBGH3kb+VE9I3A6ThCBscevIWq7tU
AYsWfLunNhrtn34nqjOmqmH1PgJcq61zENcev5DY32gc/W4t6suWrWzWXyd0lEOC
RAzelpz1I8BSEYeJtot1i8xTuBwtVf+RvPV1/r/AcAYfSu630vRYLdhLrX/HV1Z9
2+/Nr4Dan7QqpdBVIvx8wgf2nvycPgJhssmD7WpB8f1V4w7UaW+1YN5nno63/5wB
UT0mYXnJv2AUaiAA7w4vzwhROv0trIscSzRBtVCxKHg6PFHa/7IUOFfo+yKSWqpu
QTjpLwIyY5UP+CiWWYikHTJRl5svc2wExfgU8OmljZz11/npJZmx9AkCM/eIUp9w
ftIr5C5Y5qKOkwPTSLfGI89DsDpSwU3XkbCLoVzxNBz6eWwTe4qr2MoatrZN+tU1
8QG+a4oHx86saUqsz20HYyaECmOex8yf/eLNvZzq+A57YqhQEhpB1TD5Ac99U5W9
AfHZ9gXWhxjrHtP8OUuynuEHuM/+QA5tjnO4kp6G3lkDBWLanhN6xSUPkpbDKgeF
tGXYMTFQYh/MMJ7AWrxzgXk1J9czMDs7FuAszytbWAO4YT1r+B9bYKPPtRxX1T81
bk4dQ8+OoNzchl9I9iIVDXJYniZDiQ4vRYCTU7Ta0Gy8vNQDRQ3X6PyBMPHw+MCT
DB1pIUW/gYbUDH7cMdq8IkotFbSxemEa525/X1VzDjazwe3vJv2jn+okToLWZSLI
5rFkY1xITTZ57rEXJESKNVcNBTb5UidUBI6u5KpC5v73HUVCM7P5Sf/BDFWRE3ii
0X0VwCdXWatpqV8A0GjREH/Xwuh7Xf2dUHcPxjkrH55JNp1xYMDP49FmdKyjv3Z1
YOZzZYMqg9X2TtNXFfAzi//Y9fzM+OTe2vFDX1k/BC3Z0Pw/bIEdjGBAuRaWhfCE
gKtAA+/dBYvEQ9t5Ldj8qx03orOQWD9DzDok1DhzP8tGj3L635dOb/qGibiH0JGY
h4yRv6dNWNbAjuEDv9XBDG6Sj1lAgqG2vGiogNgi4m4JAJNduHnWwAjSy5iM+UuW
2u00qv5M/aMOsFRxqwRuBNYQyxShVG7n4AUkMDlFdTFXWsWJWrB+MBDcOKxye4nf
nChkOM4HpXNhl2akCoMmsw5idhdtpOSfZ6G6os/NP8fo6/bP18rxcVO4TCe+FM1i
WUUikp4b9jHsO0Co6iAbFtVJVRtQdQngvMIUfUnYNr3ReZEx2yezVex4ppltzZhi
Mmvu9sBfG8jda3e6bDwduurgVDXa4rRKWYyavGwz70o9/qAeGtI7JNCgt5KMYhvk
eqY4kPY9uCDUDRtEUrW9YA6AflJ6/w4vNxu5OUUdcpo6IuMrtCaO3TRoYwlag2Nx
plBbQo2Y6JY1+kVuQaMWoOEXEye1dE0hAAStPzLjtovOh5ZnpXS3CN4y6UrgqCfu
ofDLMLzUTNX1COLK/px92+AZVt2kxhKeVBOYcO1/Nm7y/sB/q9K44ZKe/DmJtk2p
0wvdDUTtlMX116muSAFdfMz0KMsObecuTTVo9Gnt+4zjpujFiuJXI8jnPHExHUv1
O9U4EydH9fOc5s3UKDan1Dw6yFW8LYqLojcHxN0dCBIbN279IpON4wZimCBXXxyH
5L/qDBleZt09sS9OZNr56+OjW+yt8xum6lkPI7e7+l5WOyiku1IhmYaHkPs+UxeH
GXDeUEOW5N7BdzgQ4rEklGMBO1b9w5lDImzt1Jl1cspaJ/GhwXhkfGtuD4iKUCRE
a4bna538HvW/ED4cLcemjYCCT4Fp9OQC08qRFZvaYRCVRmgMfjK6rk8HCIDeR3sD
emp9DHEplZPeMQfco6kKucWUjb2PiV/iFXAtQhV3nMVZCyIX7YGa9vZsBN+tg2Jt
cb9hAhQkb7AA6RTzR1JT0F/Uh5IgsJ4DCWcKD/ZeaZOVJdVbTJBU4r65Xmgjz4dV
I72MYvtLFn/RbqlI620ZLUg89a9laYbMT/96oRzn11JPmNweU7RmNf97HTq/e/JS
qGUu3qrtGEtY9/OzBhliUCWs4dW169X7vUMHguEcpq65Ko6wAj1051qmPuJDGAYQ
j69ta2kWepgTQC9aBfJllbgZt50eN3TCFa9K1T/L1Vb7kfyeZ+Z2YrUsVjVo30ox
o5V6i8xFSR9PYUZ0z1mn1e1avErpC11KycOVL4j+MGrvySRFvrF2gORKnkWjtne+
chXrJa2YQEHXNuCK5tIfAO5u7U+dhDW0CzSOgp8JjCkr5h4cQ21r5bQykQ8yohYF
0uvOoOwWH7MqdgyVq2Moj218d+3QCCXVbhYPt3U/Q7Uugw9h579GPPncldNElTgb
52Hurfr4ktUeoxKcPtXnWErevte+wgTEFpAeDzW+CcFDr3MdBZMVZRgSIQ6q3K0a
M0+OcjEJWO4zuaa2A0N1dkFLoJuj85bj7mpulZAw+zwb5FHe5jXjwwXFQdGXtKPq
LmoE8/yKuJRow25k2izDoq3vvnN7wBkODMtepN5gKL5D9w0LOglK+G/ILHHk4xoG
GyLnSvfZiuI0RqeAkiv/oI7n4pIpKOi+KAk15ytbhXXxh18v7UDbMEJ0W2JzyuJf
56VxSwJhgZ4rEn15oa1yr4chgwcmuP7TicPy3JElK3LiIInI0jo680V3cxyJ4fxe
TqQb9s7O4Vx+ET4TvecSK4TbULO7Acipm451qokVIIMLlmth6tmNkRcbov1Xucof
yMu9QJbPe5l5W24oLEZUnraAWSg+c8fdNsEnQxrKIhZ78dHNPzwJxXJZZreaqbkm
aqQDEPVelZRbPjoGUtWme/fbavKWATW3yKQyOSHgsn2jOcdwbiMNkzLiY/iMjYyR
ktVV1iqRwNQT/p8wrZhf/pOya39G5emhDQtIiUf619Yu64DDhjELjKydr8jPM1H4
jI8h5FFCpUfkFTuTc1jb5IyktkaqyQb9TRXhG0urSu973KATPtLKVc1iBQsR7jXX
3shIbz+bKkYaAiPCuDTD3j+Mcv2d3qo+r1Bczs1lhxceEAa1HQUzz9VNwV8LxhJm
IbLyyC5ry5fihbCr5UUEjOeG7grAsAslODAaf7Sc7sam8qsm94nY0VSkBEALccD4
UgY+NegzlOSmpbACF3gsVUwSnTSbQPLno0cpccQe+RKHIgUEhB4cFLGqt8t5LvjL
pgQnsXsrJ1UZa16fQLZb4Rf4+pp1vKKwVu8t9iKGQ17IN8OUq7suEGIlWCk0I672
DlRCqnj+ZRQPW98QzbGoUuljPni0e2Bhz0Wb+TyejygtxN4p1J1uTIUIOLYgm092
oTrEv+Bi3rKFpcBW0cOk5AW3T5J+erN8i35yWOZeNZhhsgrMKN9l1gBD34MUowdg
HEfBQltWO/AnhFeEWNuiT/zgFuJJEVfJ92n/M2OQwgp0+qYKi5zlAq/BYAF8mg+N
3hpnpifki6EwlQ8lOYVvzZiIel89Y0Ac8PCmCA9UtDYN/U/LSZOmdOORdUvu7RMN
O/hglNdbpIZXLjPC0cxz+UMD3GD365sohCOo0DJNxn2ClglXmusZ5xNzn/kIvD02
d7NTO+rnN30lKodxiVWH2Bnwlv2Z/2wGgps37pWt/XZn4lAfD+DTfZlkB4LnYBrb
bVxZSL51F3pohFrU8K8bzZDUqUvjaSNg+2TRZ8ZKus9kLtuwLSdG6BXG4ayNzKR7
jSuLL9svN3XR6vXjinu73PE6xd/kOD5tT7cxzQzCPLx+ZjAr68UJyAtYulQPNAjU
HGP1fD99vjTvvDXtwwT3BXbOAsUdk2xgGA2rn+NMlnff1P38I8xpyJQVYWqhcGlb
V4v4kbWFd1S1No4e9BNPsBYf5Yi2r1RhwXvc2RNqb072Lbit56Lonshalu+wsisq
cpOeKeX04LdnrpCMWwv33niB+AVK66jgeO7dX/rzIbaZR4ILaSItJX2JjBVd7Xzu
XPCaKFnXDnDqzStCM0/smoDs6sT5MOlSY4loubnvC7riTO90XsRWxz51iCUNoP1B
MVKHV9sg5BTjKs6/ZcnZAxRDhcWmTXYzEqKUtwgGUnYXaprI6YVT/tqdN+84d7E8
qR+ZPP+PR9JJc8fARBT2+BdI5rx7zO3+gFa+i3XZr4sxPeaumNWOg48odDoajdRZ
QlMtPeILcWT73CTbGzAiYTpIEYKHmd2IT5nIWTI1/V1wfDXp82iGfRd43aVTib8h
78crzUp5rhYW5EkU2lBSJasIk+mTtRATJiM/qAt1TTKtBHpraVQuKdiG7tSllMTv
iC2wsszvFTcso5fTtD9TCvmsDgZ+u6O/4hLC/hVh6eQp29e2E7Ccl5p+1vnA3olZ
uCuiS0ly10XPjFbFOwU6WM1jdpTQZauOBq3o/+IvBuXBDKJbfoSr5bD8VYHjS1jQ
fDWHcszx6tXJhD5xCtzPyvp/K0J7VwEHjpo06/5IFkYXcs2Kc1hQkgBMT7RWz1Wl
3VPPyAdhLRdygx/OK97yuBevVUlG9I4vjIeWXXoBIHOnC+UjbSCld3+tDCk47g7A
iXPITpbjgrenYEDBAgKozd76Z6wqvm52JjBswonULyIwjB+4H0fYdSSpT4KR6+Gg
Bp17uR13rLR+K7uQHhhivoj2bgV7Kl+8sAbQqgu0/0dJ/G77Cxkeaq7EfbDVYNI4
X13sTYO1YO9YFi4R+0QK+2PDDDwkr6Bhhsb9OnqWMBtpKK1bvyM3Vd13rX9rCpgK
DIUFXzxD65y8HgJbRamoR9B6TEGm02rGTxhC0hd977p1WrRYDxEajww2usAnkM7C
4mTAGFvJBLZTYNVZkrP5pF0U0H8QMnpd0j6z1j2OQ/sF+is/uK5Ikwxlzy6lXQgX
coj1FVp3M3PgIWYi6ovTWAx35PnNoHEDSQBDsSv37TnOK3wmOyhDsRkff5nV8cUP
aj8NRUblNQ/fA8BJtADDL7kOHfUzrla2O5OvhZXvBr0HqFHFjj/JitNv0WNJQ5ZN
5WC9//WGv1go3nAW+kGqE11P6w4kDDPOPNNBK81FqNjZi0CUMGRCPWaQxV/G+YjU
untZ6ZM/c7FM9hDe2EMKu3+eIizOJgczcUHo3G+CN3kRI6sXYz3AKY6V+eIt0J20
1JJJ43PUzPUzWmCa5p9FfFYU6YVBys9thrJOljIkkQHVmlne0WWXW/asqDwn/JH8
MvUxKlUGHLCxS+GrzW+dY1lkEk5KHRQoYiIvcaSZB5SS6l8ZUWHy1k/EAMMXOas7
5UZPmPSnokUFtig2qjaC1C9SaTRwFQSvRZpRWGrfN/5cGX9Fs0cvOx4O03Q8mwgL
TEy91xIJTz5G5aTn0d+D3KJS6UZDnc0KOXdpza82pXYygGBcBHyGPElT8Xm8AVlX
OMbq0Jhpbvl5wbPYqpvMpAracgRBXFYtvsZ/6G3KVRC/sxlgfSwhvi53QZLhSKcv
WpwOZAe2OZ+1yYGNDlpABv/fjxRNTdoskB66pyMIegB3rhtMtfnz7jf9aqsDP5Ap
5354p6q8OqgkDL4tR4Fh/QSr7sA6ORGoonX3FQEphptfeB06TG2hhmdMH14BKbsv
KO3I9HvjiGzX4/ps3b04sIYB3hAal22ZNKbU1D3RrZ9R91OLkWAmgRCIji9FO+lM
fkbVsjGuxdTx0STlrIgWldpd72Yi1bVH9FZDVBT2ywBQBGN+cA2m+3Ns+PYoAXhP
NhhjKc4Kp0l1vFHRC4YmLCfLWerWer6j1D0YVgovpnH3z4ks/067/zvsv06VOm3J
VBs5LmHsImTfRJXNQTgt+vsEZuy3dRqM8mkAVT1DpbVo7C3RGP1ehRphgYC+NEDt
DJ3cD9EpxE95KWUb16Y68eAclruN3+3RaCUpuBA7NwWUUgTIQW/MMLKlVBtxhkq4
P5QWb7W2Kp0pvbowBANruvPM04ciVdOa9yBobep06FsjmsUc4qBtqOUa3/i/umbq
sOqx9MZ4do82Bfb0TaK5Ug7x/rYgKub8EKKM/TPl2Eks177SMcFr5XefDlnWzJGw
5OEnZZE1JSvgweBOWlEU2WLApM8HFbHRj1B9cbndZCaf6qR/m+GkT/W8cvsY19hO
d8M/evWCOHP1tUJ1nUN17rsdMRMwEhQMp9QZREuqT/OAnv1IGNbDxtPIkfFWMDeJ
NZrVZpBsfgGK3UshAecIjeqC1bC+vN7iSIy2lKxKwMe9wvsbiEFHr6NPZ4iZ09em
h6+WeMav/Et4kJz8fehtUAXesL1blDlQwPHSP8Lf1gU/N5uOfl9vFAaZsVa8npo6
ZU8ADAKQn7V4MOBByq4dX4/vITrotLIzurRekZYkjbjKFV4ZgB5Agc6/PNbYaMK4
C/YpQrgym17A6e+dNqZNsQ2738DwmgepKmLZ2warXDLOb1icDnEz2M45GdnvTJ1X
9R17OZELa7AsqvREZkC3F9VULddTcPdajAL7S+4yUDiazT4mYRGOAbUniNQdqRZt
xI5jKDQk6thpRPoqS1TJKdmivUda3WUWNNRKyInxuQ/lvT2ZOHRRomlM8zYd0iWa
JALPhh6EuTUtcJGBJ1ZRy/yZWlo652wbEMIvjRLA9cySuXq8F5OGkFtahKQ8jjuu
tdMOujhQtkm9WveH+NoqVvdnL0rd/2mbvG3nX9odJshN9kdW7o8Z71pwDKyzzNr4
jNJWr292bhr+/Pnpk2YTPBOojTyZkFmAXHrsZ1PKF5Sgd7yuZBlJggc/bZF/3jBL
88PUPSwowE21NVH8MXKx9qey+yHM5pkpsERmrJ3AkLNhArq3hdN/gI4tHtoPgkvs
uAeg8+Su+bCh2smsBfJfCmgwnfNNR/WS+ptXOXAXN8ddJDZvQh1voROOcRtsV6j9
bkmmx32do4h+ejTbt538Aw9Ltdd3IqAk6H7zL32Yx6sJtfh5Ifv8gnQ5SAJmLi3d
XXI6tMMqkFCYtqNrBmNidjW4zJYOzcynFt7lMn2R/kNWrQP9lnNDnfq6d1Sc9ULA
ZIM1FNSOzNjpo6EFVbG8WkryY1dAWqjO0U0qZh/E6HrZWviq49OzlR11Nnr0+Mnl
DLutrF99vf6QtQmDVgxY9O9ATOy7DRty6z23LuJFKPbfRp2bBtEkNGkB5xbVs8Yq
tNxphlZjTNyX+iOYN/IjegXx/MqsG0omKPsl0gWBlIsLl6gMavPegkmwml5E4fMx
arysC9S6u3nf4MvbJx56TpFkFvM7bcqFFCe0dIW5VkgcTvDBDMgsv9OLeRL7r7hS
TgxQ8GI5JRTRbwzFilhzfyNkpkSySFCZHkptdK4jw15jezx5GbF4pYzQ+wkbAx0B
NP4/r7Px3ZA7zTGbp6rkEnFYgfuUsG2XFFIVlDRhECClPXBGatLBVGhMpKnGaZBN
cZpEhRzLwIOGbktr9zt7EWdNkFuai5rNePhga9seIsDhFJfcYwb1xdiklc6PPfjj
y4PE6p0HXZ9jXf+/+tHpbxYk6OQcdfNyj708OUMuvUNsWkglbbJPpmfwNMj2bkoa
YPByZd5M95c4wqrDjvVPLTpBdskEvvhSp069j43inqdtwKfz7p9qL1isWZeOVcu3
5F61AgJAvPrEJ+SPg7rPy7EL5bD71JoPcqL4TsDrhXYWtY8H9wXha+ASaNusw+zK
kX88LB2Esc4jbR6LzkEbN4SUuYVVhpSqyTqWQIktrowV9xskA5Rwd0SuUqM55zNa
nmYvsa6aUcqyJGrEhEJCbkmqjh7Li1XpQnslr+VrivuEXQquTgXkjsMh2Dbg3DP1
XYftIpLSGJyuCF5CoIeSaBVRKm7G0LqB3vgLTdN7PAz7mu+VpUOZBZtBEp7nrF8f
qTHdZwlKIrnbcudGSpZPmCYqTZbiVbwlxWep0nK6jFfmdnLdl0ILexg3xLgh6Djg
D01IC9p65qQGGhcCZ/+6BDs62woXIKXxsiFkR5kf1nHFxiaLz45nydbDIJ6/TDiW
nE6DcwGUyG7S+tk11raOq9MFae3BiyPZ1m0P6Czsxx/MojxhjQPXnoL4e88gZrgJ
SY48ERQJa+cuvtO1rHejUkm3UMAQIaNx/UaeXL6MEMZ7ZzeLJQZFspPNUt3fSoAM
7rjZcBnZzYSe+kPXQsgHTJC34AH/ppHx7hPswvn43v2lX5W3l1nIj/IQThdJsEPS
jS4dhIJbiTk/rbo9njtmOZz3UP0INFEq7K5B3SmHwfW6An1rFKfDktqm4J51coJZ
jaOJqoMGXfSvDMZxCZgkTEhbL0CASl5sxbjBQulq8FR3m1mUQ/BhTXjZ6LhsdpUz
nW3wFlNNIilVwyElwoue42JXMMJZUbGNchB6IAQ5U/0TYwV9ifo3pURZXwvWUYvP
fkxVcc8soSpDHGyMhNoLeMXI5idbnxzLcRKeguJvMCeSTIizC2xOBFIEdFIWCv34
j8XDk/tUaRREC7fVgShQej3KvmHY1wzIq6meTV0GKra18iyi/FX7k4du6TXNhvBv
ZI9DWV1KCFcz+GA0uToaFkWrSMJo7/7nvSE3KarHBnao4Fz7ezzHbf3jHbmNAw7q
rtQ1bWtF0h78dy4I9WiIZ2/lVlvIrtYRlH3kd4IzulnGmBuRVZRH6TjODBSmm5d3
zcD+8CCCMc4apYLD7MtY+IyWlYB6gLxwUR4mogxftm+eGe1PHFSu4tR2MDbSmX1S
W+luEK73jElOW2Eqcv5LlKGIvjfuNyMG//Sj99De8TfFxVnYcJ1Towkfv6f0+sdG
a//hU+Yy5ICNuOUiBJxNKGHaxbeB+IkUwQ4X7ba/tckvzSOp/4ThPGfGum/bRWM8
0YVKzYy+JLK1AS530bNdFcdXmi7Vd7apC7G1VeKofCDZ5LDTV5gIl2mNbOBOLVvU
GybQwHD5uUFi+hrn7njfhyk9w0J4CNSCLSkzIhBGQgPiqUp64p+13yxu9DeQgdG5
5K76/AZ6M1Kv5CWZJOW6Vgt+ZXcsp08M57rvopic2NdD+o6Dja93x0+hwj8eOcA/
3iJirfPtN6yDAxjn8KX1eoIJreYYa3TYOxwCSf9pUhcfKD7S8m/6ybhq5cYm6E5A
4VdCGtn8kEljRWBbCFsurTeRwcAlQaQFHsWhSbp7vp8zGlGIOwx8XWGZQnafTJFl
KJRO+1kfr81C3VnkXVcfSwRueLn+hlo7vJdxaBDzS7v1WPhU2fY7imwT9gaOupxQ
TCjK8cTC8Oj7czID9toXYduXc3ZClsSjzdO7HjTRWheZ0KKMM0cd5yOA6LzDOKQ6
5qmDPepiVG+JwW/B2V1FePlfTEHau7ACftIVQXo3HKBf4kaRmcjuxc/J226SHd9v
r/znGdirzrk3sqlgMHY1wOpH3Bn66Je4xpVIX+TovkAi4LMOYgfTPHNzaYGOdHIf
y480e+0cs9KE37lBpAFNQCVvyPYpJ2JIKSEBhB5Ux9W8bcEJ5iiiNr1ntLUMZYOl
zem67QkQ5dCMoBxm389tFbFajCI5mfSslbO6jU83cr1FDZaMGoAvsqQ8oF5vNuQu
Se8M8BgDnBaVaZ+CGk9K8vO/btoV3xXvcPLaemB45C0e+CLMQo03SxQd1eL4CB44
Iiv65zyJaD9cjlNyNvp9CKcxbj6n9dMl7Vzd/gtQj5/8gznmJBJrgexx/N2Hntwr
cL506LofB6YQFalE2zkDnSYf4U4cbjvpA9kyqj9Q7eS/ya7dwBGg1be0+C1XxQs2
h/pjR1Nf9+Hk8YoSXlh/bBDYqK06hck9FCLECF8Rjg4CanlLJu/ljJ2yN/zw1wgf
qliC76w48fusbCW6ySKx+6y6ek0nMkzmb61r0db4pMTYY/AFMdbwTl4o8ec6+CYY
Z7rUSQlkbGC+rEeTaMHQJ+GSX7RtvVZP0Y+Iy3tO7cbgQ5ZZytP5ZQKen93YSplD
fu8l6uNTSKk6TB6fjKVbr9ZrxU3TIlh5SEJV18FW84ZHeYxzvmLElJWPSNic0p5Q
rClJZYSUMhs6h/eMi0uule7Homf04Scv4kQJPHbAteLKzq+1AzwboBWRcEGgsv99
YsZoat459vsQOpAIiI7nQMxUSREildvH6jzOunTeX/cqXqPvdt0BQkIT8HZD6Mmw
Ew//h+lxbONONRCWDGr/WdBFMveLmGJR6GOHJQY7WPOno41iO/V/yZDObtt1hGS+
ZNTwKgvtptByXgf7VygUiJg0gFyZNgLgrFqhnJxNyXQ5pB8mMHbMkyC0maDHBMIq
u2lK7nGnDstEloW7wNc0ya63DpbG+Af+NBm+VREVGLspAPyzPiSCpnFojCl9PfS6
0sYnxlQ3kHoyMqmWqbR4GkB5/YfIIA9L9lA/if7qE550vyt+66JG33JywxtIaoRl
brGEknnE/Xb8w+utYImivTGFeQ8LJeI9KoeyIFaKWOVP8k3VpY+lwHbtUHyJOSDg
5JpVO4A3aKHApK5C2FNhh/AkOCwfRZmvdxq4s6elS7b/gqdXHLSiZcko5As9DYIw
K2n3S6vilOOPzJYisBc4YU0LWizsUFn5fYlYmBBBPn6JQ6P+4vHG5EFxfLXr2NhG
yNGsS7BncXZi5NFG8/rgrMFwp75AQgAwzGNHFwM8O02bHPgEyPCnsVzNHKFuwNkb
sCAKMM92H5YPSksjm1HRazZHP3rfLEY5P+z0D5USBixC85Uo4BIzlqqZezjPIlTB
DkRn4XTgbi6v5+Swi43u8/xDDHF6o/8vuHxT0Utl4jl35oSnZp3XKENe6wmxoepL
cAapK11pLCv+vgmR7coL//Q5TVL1E2Vcq159xRoUjeBGjSf6nQcuTbpqYbKMLtQL
JMznsic1e/Uy1JSBuB/CSwTWyCVeo419tBC9DFjOrU565TcZkffPsDaGq8bXXHUo
H4n6loRXYOUNMJkrkNuQ+ZwKtoLFtB2LBVQTiYINrfJm5suvEbhfguYlYiLhwo6n
jhlb5/+DNhJE21EQZOzOk0hPRM80ZgoFuZaSKcphZxUZSDO78NduOgXbKdW7VqxR
2LbFyexq+g9VDJUSdI7+dNFhxroAF2mrTPmLe/QKS5rnlg7Rr4hN8w5OZg9zSNHa
R2ju04tbdBf3zyl28ulBfezXnlFkTuu3jjJvf4wNMa3TyYK+U3X4x5oIUpJZyinr
RKJU/FOYRsfGzdfIAe03b22CQJhfMFh2tivFeqktnBVk/J/xSi7NpoLNW4sD+qTq
zupgBrwUFUOvvlgtgVCCabUXqf2qQXu3ZXxID5l7uoHGWLLzHEYH6JRe+HOVx/LB
/W2pKFiTOt6S3yvgNdmGKZgKcKHP9EXBmTb5OlkyxEBOAB9ue7gPpMXEl+g6G5NX
b00KpA//Iaw9pMPq9Lj2HuTos7lQd86TDy2pqWLmDmHXmQ7qGBi1WuX4VqBQaFxh
m/2/ve8p3abHH55iw3T2WinDU/pgMfvlqzLQxJRZTTtjN+Y/3NY2K788wg5r2z1K
EzjjuO51W7u/fEGq80GkSqFlhatReIudPTfvTWkiIR0LC9OHGFfQlOsvz09waC3i
y7oGeHZoyh2/T3T4lcGAraeSgDZwAfPssoyqs18og6YjaLl79npiLDkeNYZg+dal
A5u1ydcB9N5BBID58F4It0nSHdCHXi/VKUpn5XP0+XezFX10HxXmY26cj1+r6YLA
4XH5VYVVPiXcApo0/SFPIwImHXAr0kQwLj95NzL2LAUfsIuyXC7Djjr5sL+Tcp1n
27BM0uwkkHe2aNsRlxzccGX5RU+o+QtYqO4YqkKwSKmJ2HKqSczLrr28lS4hDEhC
Ts1wPHfOwBnv1M2WR07GcMg4CaVyGOfmn+/eQy3CdJAm9/EAik4T4frtwv3Mb9P7
YPTGKoaKYW0o3cTyBdMS2YkYUAy6EYmPujBh1pQRUlagJuyX+8PYb8nKc9673A54
Lpb0Oz3kUk7CSqZ33Pp/QSBBRd5f7+hKf1g3tMybdns2+OZW/V6kYZ3tI4ab5dB7
fmPVyfwlpIMzn1ji2Kukru6bSveRjiG0FEcKOR19Owc7FrpRz3pghkdlZz6NCe33
0KhdMpmRYj7nG7Fm+UKlGBRygNhIEJoKhMvjHZ+Q46fxKsUEbYA5H0anyCoiIozK
+oXlTQ7uEeOWInqS/PsYlMS/+cLdonWlwOSl4NTg8JrrlW95xWmtTyu14H9XKRXv
Mwbtwkf5PgDoMqmHtN5J+kGnIyRzCGRuxADA9/mit3sanj3FX9LV/Txp3EI05vwe
irb6U1DX4ZAnTT89rSZyHE3utEKHQwrr6UwoKtLnp7SuL2Mu2hLErZSXqP7xdn6O
xbHqjiEZzORNrqGwpKNTvREPmmisfhyU47f3cQdtqwY4xbGh/RNtxyJ3GSyYBN7W
sLmleW+DE+mi98IwbPKIkthUZOjbHh4udrytDPPSJMoSJX+nLhoj0fA7WkSXUXA3
kNb1LfwYUKSSijn9mMGHXmQF1EQ3eumFoeHjG/kwZ+MAxp0iy9dvarZ+KnPBY/9C
ytFViXQw4YDc69zLQwst51R8PdzloLsfbKi38neWCKVM+w2+urhYwkDDNHF/ftaR
Z3WAPm5nvIDYsUgelxUjicMhI46MTiyuPVIR7BK3iws4UxDVQZSksQaEp7myNgIm
JLGfM/RBQ7VmzVio2F2AHjN55hhm+R/40kOzpt4h2XLF1VPapUfiDvG1JQk7yU8G
dcjzDLHaDYeDVsayIsdFm7PLcBSYPXFo+MZUUx1ZGLN38uSXYuk0lJhrZEEVjo2w
+t6RltT4KQpFlJABkf/HnWQqEefxiOYoek/J8wUNQVQgk16PMKpYQdsFw4X7eSuf
r6daQOD4PiNc/u3vwM5R3N49v11N1r7obpa04Y0V19/p3Lxr9GU7g7YlsmdjGUAx
fGnub8eQCuNSK1iqJuK+rAEExz8Wxb3Jsz1iZZ6/72dasR3yyramGpNnW06Ile8Z
fCNDO7GSM7NAwMGwT0jsTX2yNIfTvSluf2O9lE20S3Dl+2LbxMGubjhSdKIAjEb0
+P0he0onquh7B0NnljuXFS79Nd4uOyoZy91BUc5HxlTE05th94riX7GTScIWRQF3
Vf63PNxlnmMbkQDodpY6I2r7O/FMN8gWTsqmOf5EKWIgBWDK3Zg7QSc0vF/vHFTw
avI2W7is4xLyT1woN3o5/YO7yFQaOKyYBLhOyQz55FrLlubhtmfq2VyOSupBEgWm
vu2CnARFFXwFu5Y6dOxDbfNAquhUoNJjo/FtFFCur++bDN240veUuC0AN5L7T1mS
A5Cm28OzcVJZRqT8Uz83wJREBNhfO0K+F8euR5VT3/AUfgHhJ5yswg3vLk2CCJyc
3yfZyIc7Qg9kSZkPXNDBK8vDxmjH75Ru5I83xWNiaZekI/FgwaNiq2Rp7fRQT8J4
ME3d9eC2IDFr8GIFyrlVZocNS3UVOIUijKsE8c+uspsF0JCEGZenyuQyGAnbSVZh
4jP7Is6Qoi3GEmdMYNoTYkqG6rvMDfWpK83JueezO3SnE6UAgseYAM2VdyFpdjbQ
NUocql8ORuZXlbJXVf8nfwr4csLnWrSqvz6HqzM28ASjpQ+dDRHzp3bNe/lyHNf3
nhcNhFkMdfCWVbRoOP+BWDbXUKnQbdR12XDp+u8o67jotGF8iXcSt2k3mkG54Xoi
7Y31O9HqXMSTf2ryaHUmyEQBW7O0cP0qCVQmzvuUMblCuJyUMn9TUmVE1WwQXE5e
sdJTkObpOxmQPYXowfHLoh3R6GKVXFUix8WGuXLD5ybptBhRJAAdgrCMQePJ2Xtz
WEOBpo1rAtYDDOYUxOHvjyz1uMFh+60WiSQOTwk5ph0aTlffBusYuAuEYWDlZu/c
PYxBxxaJiWYOpGJ4iQZTQR56uM26g8H/9eXIXQOyDX6bvTAnG6wwvMOSsaViv0Wx
Gm/f3m0Idl9yAPeopdjtD3O7QwacPdWHh/UiL7aj+/gr5dx3BIE1+uodCY+zyZIM
td1x30OL4UjjTHgfKwWYXMEld7OyL2j8KoqMcKpMy90NJbem2GNGaNaPw2ATOGzP
yuK641k8i1aszw0HKHLBIYplestnFrASm1W6tgsr+xgHRUZjthj0/MJX9/5NmyzZ
q6xxDssjrQ3x5iZlA+2Uy1NT86ZLYz/tJsQYnCHRTLkEtk9jwkoPm3TFkx/+QEQz
QaCuZm9SFqY1zhwZnxI0PszqbdhYyoLV+VOcBvXzvycN8Ar6KqWbj+z3PlnZKrs6
gP+3V8m18exoqS49jG70NQ8pybC9JQR3RKb3hYXMUeD394ZKHLH+d7uv5oV7+oay
iwu8nv/8aLcboywnxxh/UaNbzldNTjcwJlkWD7fTvmRGx5I26/SbZxOgku7nAOF7
+n13Ylk5lAOG2FswzzVY1F2CAVJLssCEtti4/bzIvgX6ItF1Qg7vIvzH9+RnxHn3
op4FNpY9qKV/OrtPJBBkC+sh2HxZxo/WPUD89wZNMRMoeLCzY/gfGb44+jUxuH1o
JrC+9nAtzfHIglHbkpWps29FBDVgfRMRu2AWmEyJ4582sTRFr1iy/fIymoZhNS0k
GX0axVGkuHA8vAinJneoZ79QdvBff50VE88ANHNZuXZ0mhKTkweyIn/zUCdKHX/E
yBpav7iTKD6VU00UBg40NAz2taDAgGxwr9SML13xpKUtiIQGTb5DYswDtvtk0YXC
WwoG4iaGlI0GZPl0ou1fTDcWgheaqTm4ZPlnS/J/wo6Z3aMwRyxN/b/RZI0NUN4z
WLxNvmBdKiqseSlI0hWrjLmSiAOUJZ0DgIQgeVu6mgEQUmUpgOFWIbcTbgFU0gab
F0ukUjb0aLlU/6HGVIoazVQ4iT6Ds3Hub3QS+9mmZuRTZHezRXChpnXA/+H4llmj
aifGrFXuxkU6UXguaM6a4gAH8GzlpcqeO9SAbmmpB9tot6EZmRoiF+WR6wiQNeGl
VNwfFspqwjeunTRvQyfzDZ1X4Fo86lQoVaUB69MDMRx1dRmPeKfekHI2w6X7EsS/
+K0c8alVzq2ozjFiap76YxcqIm95u2AXaWdwmixukN98/sVIPt5uxIDLclF2aloo
7NrMrlfurQToJXMwB5aRQkj93SojLXDN2a0fZTmo3RjbXdD+v8r3aK2RkNm0n2Kd
sppQ7iJfMDUIp2N7kZLzQiZqW1GyCphwdim/hi6qrzUc07jT3TyT8a9djCuFmpta
aVanr2EUHJ5nY2wNfkSpBBlHe2jwuuAKFGGkzY1ODFVWXyauCEg4RVd3yaE64cg1
oR9Vgpl6FfIoeXAd3GKye+1G228+h2iCs8tiwKooClD4dgBJasdCWcmSIQz5bn1Y
PmYJ31euwJyc5mGfO7bR5p8zGswWp8zJLQ5tE3F1JbjeyXtVWAr6fFXMjUYKlOTX
DMQL7wHTGewCLKz4SsuuyiN+wGBb7W3hpyXuZv3H9iEJzCQTP6cMgbflp9W9qx6H
f/SiljwCJjpk6RW3fyh4eIWtwgsoikKm3OM8v8DV9UbQY/ZKi9NqrZFW6MTXdzFg
spHDnqD8Ynm4FK/BQQbD0hIGnF8bKPzlh8C4E+zeS9j3SD+I2GTsFsAx7fxGaZ4U
g4/GyGzR6iN1++6Wl9oWR3skd+xEk2YfWlq+eLDfGQC89ubrI7V2WQoSY63F484I
wEA6IAfKcy/2+46gfuL4iKBVTLCU3pIcLraAr/bs6eyy+al7aC/WfYQPXns/vy7U
JZuEw7cvPLtHxzgDFV78VbjazP/ShLEp3vIjCd4OL941nPiSHv9aN2kLNK20Uxyb
PEl/jXi5wV2wVv0sq6dYuK6jHke1Kb7GS+oXUaJGHG0lWgnK8kJ/fWQW1hoXCgWq
KN3yNwhZfz5GGbl4drkRRdLo17wLkNoRRS/DzaiF7er9ZIpkN6zJGIUvCxQVQzQl
VGlgIqaJF9vZlFs6DELTeBjTo0jWvMsdhMqKLOMQkneVMuer2q2qnGbJycc7+J9X
0FQUX/N0NmnBqWzPgx/mQqo/1esvPXYSIaRrmj19PAuiM+abCKRUN8n0gH3d7IZL
UfRa3+fFOFkfoxiQTAEb+YARzbU/aJkXIOe9+8mgK4GC1dnZtYAIsiz4wxuqefrT
ubzX6yGZLQ7s34JCPRhVdMKKM7Svuc0GhFaO5dNHTKw0GN+fz9YiDxIzCz5f8gOT
87HUGozuxkiHPvQ1juIjfQtzuoYphQYg6Jqphf8/RGbIccnB7rR+kBRRAByCm7Zk
srqE3aPbM8IpEN3IagbPjxPJfO/HfDvTSIaqYt6MZ4gnLbPYoVPA4aJqdSCCsOwn
TXNbgd95TJxYtT+DxaIjXstnM2CdAedoVNxErEBsV32IBgGxkuu5g3kNkN5S0s1w
9VKsh+zXisdL2H0E5/t0o6PyRPUrq/eXNd6RPjAt+7ipe5Dr61DavSolhp6oZTcT
PDoFgFRsTdu/m2wGyIQiQDBZJv9cUSU2E/lX/W2Klbd3a36W/VZ6VojOv9Rk6JYo
8D7yGwsWGFa0owRZT8cO+AISqhryAveuu95R8NQ8qehiMMFrsU24iSaD4oSDlJgL
Pn4P2EG29bjGBRGl75O9lU64/+cDiK01ZAU4zEGBhp89L/X+wgP1jarDU01uM9dQ
6qOpx3C7RcVPCJEkSyt8f3u2SCjKJtivEfdSjBrs8sSOOcWXRAwsq0iJQ8Wop1vj
SXkxQvmQ3dw+pYBI2dv8PecAFYiHvfH4auurwJCRhDkFXLf9uO7BTbF6PRngg6V4
YjK83RAylhliPknPB8LyHqktAnwaQCUyoyAID3R071P4bVn8zk82x5YrvRffssxg
ZVlMcaKJThrQg8Y4nIrgDzl1tLmic8LJ+1v1ZiUrjw8HWWNaLK0nAwnfOd9S2u5y
M4P1U2Z0g1C8/E196B4G90LK0gylK7DicYz9TzAx+kuZGB6ESxOnpJJVg77vmXH4
jlKgnYjniFATC7kZ1uaDYFx9UUrH3IF9I31p2lvJgBNvKUyCoekHh46W/Nb6wfzD
kCdY8L7dirgHq936TnaFmEZjl1Tei33PTYsv097+RFHJNpD940fyyPR2VLhlPN39
ku0pdorCY473zc1X8F4ouwS9UXbRJHxVVKpoaLrki97uBWsnNKn+xtxukjPrJG48
63L4BcGfZzZMinITn5r4NausqFqBTEeOIrne6lwOBbWfCCY2Q9CLfWS+zmTFo3WL
Nd0btdZq/+NyKsb5vvdkyqB2NsjYqbRz1paOg1DyzicXhcWvuPIHPBmsYH9taLLm
ULcG/y5jhlPBwLx28s6aWjmjh9RqUIGeeoLlbctiU3HhAYgNKxs08Nl0Q8KIw4w0
TYOyNlxAbcs03vI2CHUyCNW/MEY5tPQwdhaSl4VN5o0Bn8MbjRSGqe6ievuD8wls
YV+EEB5LwPfsGHXmnpTdNXAHlbz/qU6DWPu+Jvhr9NBUIGNZdfYvhL3vUcBQ+j+/
bIeof4HrzWtoxSi9V2Pzx/tpgzuI4/l7+g+IzU9Rmx2Y9DM7Y1F2pVC0bd18eOui
zo9TnYd3tszsEumh90hobCbs5VqcmvcTupYfyKh099jGsfdiatzInbl5DdljjAyF
NadDpmCivBBrNykRZkUghFUYb3f+KKsKK6ocITygWjmndACMqItyZqq1k+dPM2ew
meduHexhFZyPOkvQ+GQqVcJvtRfZ/RAfqG3ATPW45+57jiPTN5MKYS8BTfGaKyd/
QuBghu4M2/0zvbkbh+MwqwJQFNr7lOQHLY/rdymN4PQcHls988/PpCVklg+7YI26
QI6jx5nRlsAnAiew1RSWQyKcUPshbUj3gJmcp3TJBuVYZnPLbDAYbZgxznL0bFIU
6FbMclX5VGe3dR27H3EGNtlWTV3PCYFEH/aJXstddzvU+Xk6v62lnbSVhrfr/Ib0
+KhMr4c8sLGNOcrCJ+t9gC/DJf5+lhthvRj7+Qj6cG5VwgT6a2zwjE+J9Vg43Jpb
Y19bu5KpxkVgJItTrS3OtGnYi/QRGTdjkIkanU6+Cuo7nAOqJ3RsbYJWie0SnvJz
CdBe4JBecx0pUQ259ENEquiEyJdRTfNx2OEwtJcZSS8d1gUnrlpK+9r4bOr3VA6b
0O8c/4lI5ixapaLshoclABXXHhSze93vanDp/YLbZMPMAdHL4+z4+MxRlGRSl8ms
li3NIvpVN4yqxxByW6G/IrAmdNN1pOaGqlc/dZbMWDUyHlvn/5nv3Q3iiSP3hS28
ZSlkKXhZER0em6jRFjh9K0lSh50JnmZz8iHcZkHxbL8faKpjU09WhNYQLmSoqxjJ
F3XRAaWJGb6SH8ZvkDK0pxO/TKlY+8mTs7rFoeIZqLfk0oemM7DbNb6ECtwk8P09
MstJ3rbcrhzZkfZJ39HTIw+OvivJsc2aY/fjsNtsvQGjZHemp8GqfrS3ApXMzCeJ
s8BjoMIehLrY8UfGyar/AkyhlOJkCUlE2Wg+MYxSz8dN9jF11E0UlVFVEKUsHR5u
v3LC1ijRYKpcgRHW1B/DjmQdiw+ZSQh+XuMAX0hxQV41kZLc+9k3GQFDRu13/4RI
97u1P7X2T/VI5tq8EE/vlntNkm5vV4+QNWmJq43JE8L6Q6dYSurZVLS906ZU0lsy
UEBkY5a37F+L1MjjS7/bPpsCsASfu1K9cUBrnzbSl9kCUgWpgg/Z8wZqECBfYiTh
2eBlgOBFssRzlD+y9h98+dyT2bNByx6GIeb1eUr0HPzH8nDLAw1dkV1+qwdTTtHV
9M8x8Y74ca03m6lO26Qsrie81Sht/bo22pW7FXuQ/YdAONEKhieZuOicvAQ6rV+Z
5mZdyV2kMAW/BhG6mZDKWyUyhiJ2mmcM12upRdRXv4HMBiNEIusXWirAbmmGzGA7
89y1l5jf7JFJQT0NznFI3xJsne9VVj3sJBRRvtAUJ6+tFBjuEsSIu9t9/VywJa4W
0OsGYwBjZjGyci/NnKFA8/4HQs3CEtex6NW0oFOZ5pzLpN7rlied4aIQOUE6dTLx
NZuY/GIdMc5t4dOGCIGoQf81R9XBy5d/QOhSkOo5aYOGZZI/8yDK6L+1YE2wNbo5
3SpvjqL+995tbg6zJt6AlKDqj1X7V2UCJC3NNubVKSCTxIWZ7e1AG5mGKZI/A8b4
h5WmJ/6UOamW70TaGx6nAcdf1a0U7GXGQRXBeEwt7/ZbALsVEyffhvVueBMzM8cM
MsJlLkL2mafDTnj8YBNQQ6KxKNZ/uw+9DFvM2ilz0Q6Y2Uy+I2wkQEv7vQgdF8Ug
wtoqh9a6gYgSpNofFlU5/GxU2EdyT+6Q+XXutb48CaEAVNQEeLL5ITQ8I7bUa/Jr
ijBfgTEu+/ZTfv9eTOd4Sl6febMmeWAUEZlxT3Prf7A4udSjsDqix4u5KM/ofSFY
DSE4fNVvSqjbbr9/kYQf2+PSSqKAKzBioCqFe/3atm+ijcylilJtqLDyi0kq4gOq
qpR8p+h1z6OYhXoqMQx+eQV0SCXQ3moV9r0v+8gTBGRRuARPoyJpnSLrLtTByDXG
TwaPlbcOoSVpJiMYfc+Ydi6T/3qZuKDvWoXFrNPEpmFYla7tXd4BlCS10olO6IjJ
gYNaaEIgPcpdf1R4kVNIDQKJ79kFsLZBMhiKUTVCHuO7ThCocAwBgmQGGW7tkVSg
2BCoscAHVi5qSJveocUYAz/dcP9YrIIEdynTO6EB93ofxZ1P65+5mBGGHx/NNhbJ
bVMH8FaUl7li7IACx3GKGz+5cxVi780sggabmMv8W6n77k3lFrSKaPeYL09po+nl
97snNvx5bUGJeJ9NSDwX+O9uCI0afziXIXexj7jhlxiln4skeBswCkbg/bljYTy+
RjDaq70bFOtvYazkIovWxH8dmv3bHn3ZmxP89pgabHW+OhfeViLgmWzDJ+Zk8VCR
G2kJmAxqmunWoNzyVb0MTUBNM2sWWKYp6hDY2lJKL9VG8kaJuFq6bzZ6pXWqpGk/
k262R77B8RdXmnHLNvI7lrod5wyAyz4vKSpmopc8HOMUGCXx4NTc8xm8lolp3c7m
jpGrLENZuT+3UTwdN99UaKLrssNfYQO+XNWW7NYbGB7Y0GsRyCPc3vpXvMXde0RV
INxUfTeRzOIopUVg1SQrv3hAECVJ353Gc0SaEOmBW0I+CJ9iuKsEBnwL+d1UPGUr
VSdjgFwRXLEEzySaCQeFXms+H98LmmmCSj3q8O9NkyMclqFDeyzhMOisRXmN3TG3
e7gw99psRcfR5jtWk7O4me1ypxXtYVq5f9QaMwdKWQ1kxqaRmbATX7tIwJO5jfNS
GrX3xJauCIW//OAl29vk+zuOShugVJFnJ+fejUefx3wM/qqtwAknri5yIgpenIGN
Dl4u4F3JFyjraSgSAd0BES++OeNObFUX9KUheYIeCMRmDYfR3+wK9VlUQITqm88w
E6GfnQoD76y5bJZ1Y18E0TEsGNaegJ4LZIGFMSAfnRFjW8Sz26F/RcL33K7R3Plx
MJIrMMIOIU84aOgovhc/3vA2t1ghmIoRsH4o2G8nC+dNseN2IWyj70nuOn8tU5bg
yrNXYUjkoP6qVj9WTkOZvSC/Ztu16YcYSSS9RxaFjzRtP1mpy0f2sOt/ld0DkJEX
4ZBZQ4T2YV7b7WlvCsyvEg3TyBMp/t5MsF99C+itl620WeOCfnNSHrHpgmfYAz45
SyMQZ2VoUi+/+4y34HtamVByM625axcf8/3GE247RGFd4n1BDdrkNzqNXryDO/Ii
6Rj1G1bOMhqIY6T0UQ5P3bcReAyvHGW1RqgsuWACacrSDEzfVuKgq+f5y0UaeLdz
tnst1ogcDEFt1YQEVSL5nkMgXoxdubJs/PkPNjpfk8KeV5O7Kn9t0EYw+8ereLLh
fDhelEk6/FhY0bEcN3V894WIElntcbSgBa4sQbWBZ0WLUPmoWDnWhhW3x3SeJlUF
37+63YRqzSBGaWakGKucJrWebUaI/qaBochwK8hRktcqPRQODpaZx1s+mDPjMRQR
PFgGP+VF5jgPuj4uc7aIHeRjFlgFjW3r6/iRUft85dYaJ4c684YEtTz/HThQlRiK
Y4CFij0oszpS2b7d7pOnafsBQqahmj4zceOZSEQAVKmWMEOJO6zztazDrmJLtZmG
II9M6YdcAYZtMoTXCZJedUs6YzGxD/emvxZnybXbZa4xCZFextX2N8hJO90ka+ch
VDlPvdVDmzLdRxD1qyshSTYfxRm23gnForplkLGbRUTWMPjS7MOd9HmHOYjjLkSm
cGKAnQyq89Ecozd6YGm8LjPUenN5XLl1k+siLMrAK7FHniSzrGXW84mPCJsOVa9W
SInrLmt59L2Tl8wmlukuIL7AkSgmqQoZcP/FbwxhE68x1aRQYZSsKVgEorYQMjdg
5qU/H4P7MmBUt9sbqCCOSxgOOXeB5BD2ZHHzSH5PzCFg9X8jFs5R+AXEMoRIRI69
dZcSK8/CUbTSIc6yP6Z9mKtmMMif/cwFyhsm3xR/PYTIvNaWgMijZLo/1dFR5YOL
SxeVYjrUs1FsTi5oBSzyIpze+csL5AiCeoq8Vl/UYlEyzsT3tZUmm4PX3rjXnCNU
S9yboC8sap+7kd4LK/mVQ/FyPFjUWtZlZnbTnnf6iWLus/wXC7PEPxUEMNoSRjtM
7PE5BIHhN9aM/hZ1xwNy4Hea7pwxDXP6olFxNJQibMOxQz+N0dQW4NAgIi1nxMrB
o9/iq+kj05FObL6ELzYA4hI6KRwlyLq9MVaOnt0MLzkW6lwj2fsfS7uRuNGVjv8b
37llKsk9RVlersO5jTwpwNCGs2NLqmnH25EtU4u5GGiTo0PWeGjxOwxhyLInfuGZ
th8sHeMtyRBF4VAzlGRW0ZNoz8pwwoDwNnOHQFaorFD14DJTw0ZICKM9fkJGNcEs
b7GiUfDwKzH4m04EtUllPFqtCFQuSGRbq+SO9G/pujqgKaauWvW4KyBjDxDSgLNO
Srte6o3wGgT5ueOMepmhHLv97h0vwLWv28ruOdil1n0TVYuRHgSVQNMcCDQILzj6
+spHBwHFKTs3E51MLlMwSsKx1EMmFtWN7B9dhjIdqx7Uo0gljJEGRyEPVbRD3t/z
biYvV9v6w2VrerfdLrJBPaUW0SDz2o2s5eFEKNDhpxqxfKdztGgm1JYvbZqJgGJ5
SiJrqbEI9J595fuFQyPrpF3cTwely3J+/AJztPEOJiXmqMYN+9A0ev+gifYZiSaI
F3tlntesaWqZvEg+QsYonD0epRJ7w1XPSTpyZlVH13bt+6DqHMBwMwVgJfXok1JM
yvcRNeGqX9MRm9cdj3BnmGTPAlK927R9iHcrYJXpdRNd99KrINBmxt760l6SDjmn
1KQYv8PPg04h2bwdmg0xKxoK05p/qOrwMkdRHcK0yvvmiBuB0pH2JEwIkuTOgeYK
ounCOS9lpMo9M4Lzo8pHWI+6XmEmuJ7FxeFja4zo57hVuMkFwuMgmmvG+uS4bpXS
Hh7HKOOoAMYkM9ZrcdqNtstSdsJbLL2ugoHnjOGVUeVLfg+lI+vfI+6O0IexnPnI
/vbZdzU0QjGYaQjQ8HVnKK3DgMo8mPP0pGVehrsNf8O7rCYxGprErjub3cK3fh9S
tokfi8PpQjbP71fXRZbLk8+0QFnSF7Fgf1dd0eW4NtBTuRa/kBQvgQEWODWTvLKR
rvyYo3kIyMi1FQxNteQEAB0AYYYzM8fL+/ZENC9ed4do44RtdXxYPc9EeEKs5buj
xinxnNcS8JonHx4KsTvqC/zRG6jI1w/q6oDvLdcEqlyTQ0IbM8y4H6B/7rno/Xlw
6uALAqwt3irvGOqwW9PxNXxuz7epzXiu11+TAAHqYCkTePxdV4TPIm/Ee+vns150
4Tst+Ul2oLQc5L4oUda/k+3vG5XeDrE2AdgpbCgWZqHhAp8NYtv8b8aQPWfvnA3l
zT00U3iW6h8GRKqMNrdqeb/K5acD6bFwQjDxJAphF6bhaViAgmWLT9AVBd+cq48k
lqus955kmMc8ArVmjedSa0cT8hcFs56HDE5+hm07Y91+zXuGsTUgmNdGrRjkbLKq
Ekh8FpFKImuGdZGRszJfOj9OrFHxzb/fBtqXbs6GaTYK++NHD0haoHWk/rhpieLj
jYdk5ChzFlhrYi9kFHjt4rQrK6LfF2wZiwFBM3yfBQtwFDx5KzzolYFHNWq7Asy6
WuLTOzLCCeCVXt8+SS+zOLZ+d4TphPF8fzvbe1fjd2znZiNbfwYYZYUHrXbEvTF4
xtGIgOUrhTEnAsdp3aZd4yfhHLKjjMl0NrO4+FZgZLK2h6fiqRE/x/GQApxjJ8pF
awE6ISOjUi4wEC/d9cZrAB9ORCbhOBu8GOEa9exoOvIvtZdlqkEr9i+IOA4luef0
NEOF3zuTBxhKcxBu525GMXEQdAZQ2+o66xhxSNGUkRMTkLN86qLr6BfyLWV9/B5J
CysFIVmtIYY/E0/cswR9z78CtXch1HZ27uwZfIBXFtAnYNFtwh93dnpAm4uiSvnI
VK53wMQwtQibem1x7qjSXBVldhawIrTHqzWF5Zl7U7fpFChxnHvWP6yhN9oZLv/o
6qWe+6VLNfcdyRnvtojTCF/B/ol4ftI18/4r8ONga6zKnPs+tz3xF9R/xvtFvkCx
jkrpLFHQTX59TpdczQuEPvP4AJAhVs2igSvmTrouluhz/kEE+UvOrSTwlY2BWgh4
BfTrL+aYTPG1c3fwvAS1xpmEcvd9h6EQAycp/s1n7/+KbQr/ZUcrt3Jekm13PLEE
jav0htDJPWIILXXAzVyUv0MG8n+Y6mtvP+kNMez7Vgtkm57NG0C5VfWzUoRtY2U5
3gE/8Ija2Zvm8D1nhqmrTbMWIiDnt10D67Tgqu++L9N9KMgxDXtrIWOVtkPyY9O0
9EyPOlJOXos43AyYx6OkZyUTKsiyk3Bk8FquCtEZNTYtl6D9eSasfbaKB/grho9a
kRAS8OZSQFYdwwvsh4Ap/NMyOLZeAGpoBuhxoIlelY6HVwDLzOazWgY31Kv+Lf8c
8uS+3qOqw9ZvJqDMiDPDPdbSdYfLn1Hla7EBHP6Y82e2zR7xsM4v9AWLK505boZc
X7bfraaEe5KfIZv/zcTgclsl/EumvqDuyXXO78F7qmjMzfjAW24n10XoKMyoACBS
n71S8/pjln8hGcSqrMPoPZgk6inwQ1T1E69y0otsMUonKaiQ6XzA62Dhps3B+lHh
P7Z/Z6H7uHlftHZp5g1vg+vpBiKmu0jvCBmWl0UKU1UnMkCHizoHCUVJumMgujDn
8pOzJdnnCx4Gr2lRyRs+462+J0CX/RoBEMLUAydR1A9GGKM6/DU9F28wGf/TWHCJ
3jDE1r/sYrQo7c2zNMtDKRn9IvF5qxiir60Dii/qlGpHab4bZP8rpm6UmUmTQl+4
2XnVVrmAHf4yDQ3nx4Axh/d+pWUZXpveXlCPJmUp3I5iqXIddbuDYzWiQDd2K/7f
7qAFBEWqb2QUmG/7vh27VStXzN928+l/EmoSnViuNRk/As5K+xQkh1OFStIYV5FB
zQ+XPLDb+gZKgM3qNamF3cdI3FQL1CpkqEmTxHHGKv3TABn7s3HQ/dwVNWHbFBNK
3P6GxO33P8+jcBUoW2+rAn9uWuMcQ4ymRscSK8EKmKSFFQwLI9eFAt5fPd7m27qh
55+AariG7Pr0BskrypEWIfM56rvluQ+n8PaRhaO3daG91ZG5HQIWIec6ulRP9xAO
wchfq/jTfSVytSn10b2uBFucfnzmGB80/DOC7pG4t9E5wzPjIbJS4qx0+oL7h/gw
BzRdfNJLBVl51dtcEV1kzuMrTYZQ4Ez0nIZdjYGSTjobG8OXZJSvo22Y7vMiEArk
RpMYpdb5BccQtq0QOb/CIH0KHzy/YSScM7CR7+XTfY11BVsev9po9UlNbUs+jBnu
oEl+/xER5A6tbAeLtg7sclXVxzqpilqSRALCLoTsQXnNAZGjwsAU/y/Mm4caknLH
wHKkKCaGoen5ntG3aEhoQR7nvXXkzBllihhLMbPJ1kThtWUNQFyYRfuRBefWQ+eE
PS6mrO4wlTOiUhRoevyQVfjml1ZA6cE5tClzBWWR0+JVNq7DaxxjTdsvjppN+JkI
yIDJn3sBRSkDgw2rTFkdfo3gEtga2XAJQcvrUeTpKWuI8FM0TtC0OTcdN5eneR5c
ZUxDy6VM77s81hs7qjBkQ6HvQdYnqhN0G7miJ9wDo+GXjUhp/o5F356a9sDDoIK3
0DSYyAyW9RjKxz1p0UQnkFBy7CFMws9KOyYH9PaVQBKBfl7d23caYxcBRnaSMyTf
o+PQae9hpczRVlIgntzpy5bmITKrMJzGTdaq2oiO/pW+Lj1gACITalSPjABK5MZV
2B+OtbxEJN0MpEGLVHCfFv5dC8ymNNb+M1dteRTog5T/3TVp+iU2jb7t0CzDRk4P
Nzmw2v7388eNBKQpq+g+Cc6XuhOBULYFlMaJVHkxPBOe50PVgfjEw/F3iLIwm7np
UHAEkkRmho0N1Guf0u5s1Wqz2XcKd+ezj0p5W7Uk9LPVGzy475RythhbZ5nqAKLg
legHXG4QWNJUZCp09sdJds0t61ibZcezghmrrXfqSOULDPp3mrBU/ICWayHZABBS
FfUox34RPiisfFMDI/em2XkLgtY4KFWlB5o6xaUfZ57QHzaI3fwmEHegn+bjYYyI
DAWhYJlf+fYOnD3Z6B5hCxwVB6Du1tD5wcEY8UDfgVTg9J4HFD3oZkgYjD7YSEg3
aNBjfrsIPHfN4rFLyffVSYkdzawyQk2UOKBfbkJDRsuN3sp5byDXR9Ov2XnVV0Sn
9EW/I6myEafz7QdtNYUsrKf6CK4bbK4xOnUZdb9FELubU6wyV1TaXAJI4iA7CVUK
/1KPhfvDO9uJjNmWI2QsP/3KWOGb/Ssmx+TCZpzlQysc6iuJBhH1HJIAfCjRtUqq
A2B2q1jLuP3CaSO+xXQ/eiu529GZmZcc7yaeX1li+e1zt29OZoH7Fw0XoAKlMTyi
6AXbEa90GzU/7UjNZ0dDYtDi+UICvPV2JbbO9950z+eXMiqHORmhlOVC9eQ7qJNg
CnNDDONw+Lyf2jRP8M6JfEAhr6+fdA4XQ9HOHyIdgMu5fJeMa4W59RHe68r8bwrw
2JW54SlMLExQfLOX5YDC2AQ9E82FKkRyoIccTb62P5/VXu4PlOdnU0lwGhm/3GnA
cQRsXKdxq2EO9ztOxWgB0/0YJaO1JR9wGuwQx18UbS1vAhmy8FfH9NhQAWuL4v5Y
MbDaklxWGaAG0+TShl1JPFod4qpArJ9PrCAQrgxzVJh6B2/cYCHMqGlsq9uSewpJ
02Vw7iyq+2/91DJoUC+YAVeccYAgiygwVMSITeS0H4K2LV/eCD0RrDdW3GHVBGqV
eMVWmS4f7WIbTLhjYTmYrs2FXlM9N7mQMo5xyH0ZTAcppflc75GXKy0XMScocuCm
AV1/IWyksiii5H5ZI9PHiM0secafQ0aGwBSrZX0WpLH5vti3Qai73+wwzwV0TD6E
xCFIFwlQzd2MmT6mplHYi6f+tODcf2eC+WYE7hG7HP4ch0NL/H122CtRdxVgtu4K
3PVJyQQ9+2SWBFHsfP+Rfh99v6vqiUc1pSBsotLU9qwsofj5l51ljuT60reY74vT
TB3kXtPJ2Gan8ihkt2CQ7cOqovQkRPcCZD3IHPLH5vV6W7XGLkPdO+QkcYnvo1Kq
GPbVoG/gqBJI0XZmeTo02iseQwzsIxPuk2vxDNMG5OXPExRua0MvCEF7FLt0tIDj
JdKEzCrdgHqh5D787+ig5eaFVbaq5KMC0gwWcoJzh6Q6SkJNoP0zlklYCOaz3Ue4
3BF56s6GyxIswwvpd9Jnt0LRB7gOYvRsD/EEw4B0Fys3mwsTbRLRLnQsk7swK7VZ
J5ROJvg5vDtM2yqfLysqXJxFxWbpYIRDvM8Sx1bzRg9pLKvm/l9he1HYVVqIqhA1
7RvV0cXpISARgqYEpWl7WPuGD5ijGvYHjGpjUhiIMx2d5nm3XmhaQBxpgdpJ/bBd
UYQp+FIOcSG22saaPi8npPHcXx+eUwaqayGrtCgG8aiXAESKKnj/EwuimYJp0/D2
uWkCfydTYjoTDLTd4cZUFsvEd0jLgu0MOp4GLAgwJ3BL4H6q+3fU3uY0Qj4v0bGt
shSXjWEVxzzXGWX4OfXr7XwjIbvu8Gq8QoVSexH9Gmv/WpctrgE6p1gTN4f5cmpC
eTGIKkAI41/Ud8I7SvYUEKpDncz7MQxUyi+NCM8BfvorSSh/31Tx4AteDJ2tFtBs
4dC96j4YqZyVHR5wW67tuXJuQA1SmARiCWhSQU/ulWr0rD13jRu0IN72b0pKKsDB
j/NZ4DZx8r0RP9uiMhldRpUScQMYOPMEMxVqXG2BLd4Hps/fOQxg8ZkBqlfPIc+n
qsS5qVdY7bwneDT+FQzusBJDui3GByQoxNfJ43FK0et20xB7uZSP/9xsmY46QXCy
aH86XGK5VC/tEBF1PkxmuWjZ/alzlSMjJLg6354LDTsHYquboz7h1iUhh1sITu5x
429CmCWjpIyfPE7XrsxkGmpSuH81OkvIjuronYW5T/jd/8lLv9ySK5oywDSXR28B
MdjRu20Phpbp0EtKkd/nA/voQoqLiLmj4122r8tmt/zd5izQDTEm1LE/cwkmWgzE
vahdd+7lr1gyYLcxAEqnjji3eIdEdkz6a/+b+C9hhOD8sW1H/r0CVnxdLiFPaViy
JWmoM7V4iL31cT5ImwQnIprGHtPRHzod7PyuAk8lKs+zTSt7Osqx3VbGT6agqAEe
NQ5z8lsCVAO/WcG2klRyzCbZXQoQ59YvzOshd5jVOcUF2KegdNnv5Exatafi6kvE
WDIdQhFtueAuS20vJdpLuYvj2sXMPs2+6MR7ODfgeNaeLIIHGjAkInBTvIu6MFjG
lFPIwq9SxBKZZXmkvCzPnky6isOdkbMQG6d9iQl0UGEjSpWefuBYd9DLoDPbdRI2
3N7InNQto97YP960rP0ZbwFWcgpJg31Awb0py4Sg9VnLt3DRMKNcsOdiikKkK5sG
gFnkIXYn71OblDdwEB5eMwQ4NrB7cfcAgPy8x5TFst9pC4XYIIMuiwEcM5sUPU/d
FELrGcv8zjeW09KVN53CIPk3dBe8fMBheE+dJE9bL3DHQ+20rT7M5Qh5c3AhnERE
Rig7Ue3tZuHgMHn2xp9tsjbKSTjOqjVj1fDcNkURqZ78rN+6owXIbms/fLoLDHmh
P0bIEfMFa8Pn2cFur8bV7a1CFDjBM5DkxbrCBsBJ75q4al/vVa71jhQcmwUpOqAs
/2+Wkhfi3PzHjGJt4A2ycNR3bh4rZDEO16FHrmetpmJx4axKEzpCoBpRNI3Kd+PI
CQGqf0TPVOLAbXgriG8vLSYYfRkn+B6vKpSmnkpaWjpwbJPmIayzH8WUGLIJ5oON
vhqt1Epx+TRUN3H/UiruKu7IC6n9+JWF7Xyn3CoOicg5B/Qdmxo8TFJoHSYG+mrg
26wys2yyUb6CC4Fl2giG/JmozgunJrDksVoaE4A5B+fQoibqfYZQ18DpCEwjpHTJ
rMV6wiJCilJ8DBg8O2Q4tXXyseEKmbc4xrQjQabSaH+2Ib+2Z/IapbiBeopNM8fk
JhZXRQ5ATJA22V8xkjDfffR+98Z3laoRFd8w89BFWCN8Us3FCsDB2mY+5JVXcg04
MWEe7lnjWWKm1ljaJRHmtyGAUWI3AHOKKyXccF9AaqwAdwbdRh6w6hFMTDzQujh5
hBaJ0XopN/1uA8ZfA2+2bEUsJUxIK1hsOzicP3VwH85NQuR30e5SoOv66PhUeOd9
LzgWMoG/EPsa6G/m7HjJzKh8JVaWkL/+DajIAIO9fAbcZwiHVclONbA/Ihus2pyZ
0Nt3S9NuHI1ACxfqwH8HNEmVPJqMsk85vIwgBXpOlyDcuFYz90tndC8VCVCv3LFn
aQJXNan22wMs8YyXOze9VKDS7nAmhSvp22KMt72au4ZL7rd4KAhpncOwzKA+S25t
/o/sHry+jc9sIbRGu2mA+XlGyaxD54/N59Yxh1DW70bNlO07svbE8HtILPTytiuZ
PKNdplcxul0h82ed/6X1MNkp0++VxpUrG1ciEt1oW6rPajN+jSL74HBhnLUi4fNb
gG6jKiX99ECF94oo051v/n/6ssATz6Us9nNIDsgaGLTB0BWQyP9/SLgpieOzVuwY
Wxse4l3P4u5LI2ZwG3SaGJPiDHqriensz8ouo1rJn26+BszJUe/HjvM7BTFwgKMJ
VWDNlab1U4KUbqdXIchFfYMNg5NKUsXRnMjf8PBID8/dpsYn9Wd7JzMViPNKBX2q
yi350pdwWd5ehhmLu5CjxB4aLLh7ZpLS8a7KwVAc5HUzkwnkMQnCT82PBWlT4HsX
Jvb/Rf/W82jnfkz/gS2DVBH5C+ZWaAmz+hDewrhN6zNOKg1SP6ItH/HMHAJsrbdo
2L507+SCtU/ekqvIJD/vjmoBLAch2J3IzMC8XlyD7IswGSGjpDzbzP6XAHSuj82d
ScVukIDvK26q86MA5bS60eoERUTg+uzvgQsYWNLCXNaCkwUEvlxXnEWLSmmdm/bf
o4ANiK13eWzl14C+vucRy0MY9LXGPIflmVpQ5vfzCVIHW6tBfwN4fRQyWSWKpmkR
jqfUcsTQps+O4cPunBCXXWH1EEyVM0kNNfRT4Y6PSyE9SVgdnS7it/LpvSNv3DcV
1eRjVZ15bqIxHtKPP1ke/1R4a44KWbpeAJsSMPszwi9yn0wx0k1rtAFWoQUy6rP3
Af+pRssq+DqtooZ/1z/i3t67DTxdgeYvO+4vSMczLOUxBSAbG8oJEPoKBcTe/qYg
DAgGP65b5Di6TWie18agAR2HLA+Z1mCR9IohRsu2jtxLIwS78xqwXnoaWoBseu2k
vjwbs/g2ab4as4mmy/SLNSDj5JvdufPj4Y53XSJI4RhbUJSYm6qR9BPoYh/B2cu+
62DBUEDkAwGqAWfvjKwDFQ8llZgeXJGyLNAqHB7d0b3b0+FqkEPGFnIP2q5L8UBC
oEMlSxPqzEzginWxp2hFWelBfN8Vu1m1+/4c/UeRO3TMT2+GIsLoLkl7wRobM+tv
1hzcoQDM/qJ5Xf1TTgapnvMXfDeBXvPSNAhtejWib6Hw6Rvi4zGm14nOSKxRR6yM
0YWSG+oz8rWug41lhFeYVl9BOGmWJ/ohLHYMb8l2ftbtSuuyy9rnMEjqooH5tFgL
5l3KAqbv9vALpDbeQ4AF+nkVIWxTKIshEGFkYBbEZ8OqzX2hYgF9c4cMDoSUcgaG
6l0R++GXZNoRgWHTXTcLR6CG6zS8fxuTYDbK3xMEQKd3GhdtB/gcKZwkUibxiGS4
TqJ476jvMM0oYoI2xGeWD9CW/XtnC7kWLt/Yl5WEGrvJSa/Hxks7L3z2M8ejjwIF
TCS2G78q30JXfkxPfBZYCH6MiY+YYMcjZo48UwkZNlwsmSu3InCIQLZW00KNHScx
Aq0az/39Qam7U2iqjon9x5WCJ8iVkh/+VadVLzsfxVf5mga8RWV+xLccUBssKdR7
VL04H7yGLuyYVCfAgpeDmVvDZkoAuBaAaPgcKlFHMNrcIXShyeZm1jorTW8spO8W
6ZUhiNuyxjZlnVAXJeLZrSQG5ztg4GJm0Czx5oXd74BubcZOoMuZrCHW1370hPMr
rDwzkKOGa4Ry9PY+d11UWgMEtQ7sneW9BL8kLL4CZuTArfJMRrpKFw4CZQdy71Wu
Egc1vP+EWzgoPhi2nwVmxuBY9lkdnR9elWmX4Z18C3kj+L/HyX6gzHzDIUH7I+JF
19sHRdsrweGCtIaUL11ZDGrHzUooPz/xMBJjutpQDVdHAkqn4mHFMdRVi8C9GpGv
QC/tB/XKjXSC3Kp6i/eJwr6UfLFIwRd/nJ3CkwirvJ23jSISOVlovy17icETAZCT
Ol9rp+ZhHKsUOELcZmtJMAedrOMKX144e+uxDBqvMTZzswOgfAAjmBW4kMwz/jh4
b0jTGnBWGd4PK01RNI2EZlgSXdp7BtO6j+APF0qTVWl7MXhvS58pGKaPstzB9cl5
nUqLFGQHVDtdtW+1h21mo/RaCW4Yu1+AvDWWrm9yABrqF2LFQp27J+QJybLe9SOE
S+4nH8xsFYLt2SGHzBqELDUYbaIlc2gBRcDtrVHVTSyHDIsGUvFCofCyGM00zxUy
G3kGJrOy4Dm4Tv8cuD6Sf6j07VIAgZOk3cXZtBDDs4yWMqa8S5W8eFCuawHK0Yq/
7d3OJhKHj4uiQNT6RM5ipdWMH+bhycja4GkjcDY+UisOK6LC3fVWHDctyQknJpNG
pxvn1z0gY4gumQHN4jYfo8hoUG4mJosmsyFmV1msOutKsR8QdSLcvDqu6Xcrxwxw
hatk+WC/VVU7QAV9Kno6jtVfgR5aBNMMrdC8ZKa5UHrhzAH6grsYE/E+YH/m+OiY
EcggNBBd5e9n/iUk6CDv8hBmmr6xAf+4jtOSqW+FmAg8fFeFWvH0LSnkmZ2YDYJj
W7aBixP54sru/9YBZVps32lIEwxyfBuseTu4XNpd556PQBnK5ZgE6KMUGhr2DHWO
QMJDYTeJcop6s4ZCuQfw9RUqjajb8xtVdpZ6e0iV/uYo2+gWWMlOtWQoF+qXqqe4
hL2F6WV4lrsobYyVltIzaLsvBSkF9Lg7wG04iRefU7+bEhU8HbFcEg3esGhqgM/B
TrLguQYMlU4y2fQnMN/hjkD1hNRWAjVfEmy+O67lWNl2swefQkGLpHpRaNgfY9gQ
EUZyUh2N8W8nxSVhI6Ib6IhBAer0c15X94lBwNvRHPIcjKQeCuT8uDR0/Ww+O0A9
KO9s6s3Mza4sePGUQK+7/iHk1MAcnlt/l8mjBiIe0HI69K1LF3mxdRKBTyzeXF3x
b05Nd4Z5TO7fUdTf8m5lIwkSgSbUqoe4RUkJY6sQVWl7E06Xf/8ghsrV/JFqzDAo
gNTWEd49ODW/oFSeuB1SlB+n6pwFc0/KqlKfaos2svbdfGJd57H09SMQO+ucNwdy
cqGdMnoXLr+CzPzOW66y5rm0LYXHqlKXXVf5HND7GnUwvJVlCFHOC4Gk2TQfRYfc
AFk7cFk6+EIkH3wrXkdkVUKV4LLmRsv8MJ9fCpQKNASlHEyOAbgjv+6XQlclkIGc
FK3kYw6qj5h+cocSV9PCOstn4/nL0onIO3h1K7bWYRLrKLuyc2yj6WwiIF8b2/lm
5SzQ9MgD8CaZFip74VplwDBKRK6C48JqCrTrkkMbxNwFwOALQztSZQoR9qyYxNvY
ufbte4pGC4ZrtCOmH7ArxSvCHLR4o4QWzkmnK/xb3sxl3UvMfVr4xa+n1Qh3ALp1
j5+hmgUR9hTV3yTgayV1QMNn709UPbF3WPB1/OhqCsIbRd+7YsND9HuQaWWuDtKy
Qn88AS4x+yGlo2t1wek+lqoLzGljkkyyNe5b5rF5Uv7D0M9hIjy4/IbkMtCwJnan
zo2s1yK5Gduh+WL8UyZFOdbsW6GJHVKL2/GSt6MWQVX2PzYrPg6FaGhAe67jJinF
B+wD3PPNv0kDiW2dH821WwUTSbOJAwmQWE6AULhxk+WSPuiGxm48qs9cqmQKnz6I
Mqvf0y1wVCPXPEva0ndykqq1GtjH3QM/HB73+8477JwXMdA3hMJT6Gupyojba0MV
bVKXFwaZRdKFX4LQ8F2rfk2rJ8Q8uKLCrco9uo8mgt1X9QVCDjUhvHXIA/pQBySc
1l4wkxBU5M66OdLV4pWH9OvIe3rc8v3umDUHDidZLmmhN8caXxCmHT5ul/aTJWr3
kLFCJPDAZ+LR71xewRGzdVZWzQqXQ4nbC7Xo0oXUDlcRkqyTpIYnJVf+MDHh4EXp
z0fQzMLGIS7OOCVmWGd40+akZG74GnA4MeXluDRop4Vi3T08u8dvGMp6hgeJTqJn
HRdA1bBaSFGYqmYQOiGMmkwgZ0KrOP3ABjhUivn+VQxg6/2l1zCfCvqwAoCOBREo
jXFEERifW9wmNpDf3b00y+r7tFf1u1TBnIlVApMoTCob0DT2CtQJ0JHRHk43838C
uO9UkiSS1wTLAihWeHPiq9x09dXtZErCu8n4oN736RIKnf8yeVJeZrW7PMTcur7k
dNWpyVMRvCtu776jepf6b41gMn8Yav+gjh4QK3hq1vwbDKlxdScrqOap4q7T+L0o
b8boL5w/gne/Z2NDtuXohbgAqf8jA9lSIyBIko2bUbMy7rTORMv/N+a4VKGCBQLN
8/V7E93FN+2eNrHITt6HSaKSb4MAh4vlXIrp7AAbjDXOpEFVDVQk8iz7uIDZEYSi
/cuaeRTUtTjS3bsrY+jBQpUFgc8VDU1X7SM7N3qMT6cQsZOuBYFEhpJtWudcZn1f
mwA72vvOE4mUGX+DpprzbVrVtziOzWmxI7jHT1Kc3Iqcf4HsYoWoR3xspOxqMEYB
gx/jHL+iZDaqZcgZ2IhjrURgAgZ+eAHMwhCcsqnk0JUOOYWolZBEi6JL3N/GoNu3
hkiIHsjD3j/+DQuwKWsNed7Y3MxY+RCMsXG4y8/Z1xmX++V7oIUG4dTGCVkB2uQE
vzq5FID/PJXZXRb0vwbl5C9W5K+1nLAdU3dmUjKEJhs6cwyMMGzn4/98KQS5vRIO
x9I9aCZ1inBZCANtE4WPHAVPf7FXLdwnhEOO9/T46YTn+OhVIsItDTFsXN10aRKv
GMqkpdqnxxsb6ZhGgVPvpm1SGpkkuRyGiq3q7EAyxvrNhupPzFCino68Ec8j1/Nk
SKgavgqgE2rbST0qSBKMndi8Wv+Cuzweeb7JZkAhFvHx9947e8VcZplxX7vxpt5v
NZKYh80yjtbeAXgV9ylG6gyXv0ETZpEMgIQuoX7EjyXCqsanntEoIfC5oi8+IwdS
dXmwjQZqb7IFqU9ZpeNti3mQ21wyYQJadBemvEedeqE1Z1qjD2yphNvTpQnZqURv
mxfMYtArRnOoYoCVGghmiijS5GhR5lKXQmb/vgf5TIpDTVz7t7k3mSGfHZiUGhRh
DP0GwgUjhkMNfypKBIE7qsV7ntCN+F7rtL9KZaQ3wnmoiNLax5LiS7o1OOLYwOQZ
KFzfz/uZ6zdslvTq48uq13ACOIAPb8p77BDX2XzLcfpqkjXvWTxSh+6GsTbT3vxH
tuGKlSWxY/8vlvaSiwNCHzxa/Ecoy4YQZ934gqltCPDO39djtUm5w7GuS4esXP3q
01Oh9hw/o152G+/544seO0CoGU2owe6ij4V2IA+v9ElCckTNn84JWl2PJcF78iTL
d8JYpg7qNNyz3P3vGKju6VJW5f+F8hgIYKvTKWaBqYEzi5bRVF0HGWB7NM3910jS
BGeRgFJsx6oOOu6beBioZK92iDF5JE6zpUi8gsysWTFW3bQ94d1+C4cPtfoGr6rq
4alh0cFuDdQ+yeqFo67Jh4IOSd9bkucmxIikiugDm/naiATxm/uuQ2e2dOWl124U
ffcorRelp+o7wwreoaFGmqEL6lUteuvc0NgxhadBL7iqF8aTi0E89LTpxG7XNp7Z
dCHmcrxtwEOMzWkza9gO9zgMV5We5TPcQqzc4QPaqo+qNF+SdfpyAannvZA2a0wO
15v9JJ6XmyaOm7v5t9MUkpF2hQrGd8IBtGzngjuty6gLAzZMVVJOj/iBnKyI0D6b
WI7Zyp1avde2nBCqur81TzuF3+rLs2+G/v64/pQ5TugzGn28UI/9wLzv8EfV5zBl
RWn9baETYzIxXFmTCgRQLSafI6vGYKsrsfrprq8ujsF/20gn7OJHpJa8vzU6CnPF
SK1J39dSm/3sIcpu6MkYwaFfnwP7rWjgYEhugkGiG+StuNiqbScAiTHW2TGmcJmx
Rj9TMYhABA7Sr47JjcNKmoSlcydm5tdtnDHBjr1asRe1+Z+fabfJEqfAdcSUxnUT
+txaHhsso8T6AZVUPKNIDhsOmPw7EpTnltA2MhTpqbVVchSnrVIWJr8tCE9fopTP
LMsipyAyxl1LTMm/o6sws0/O/vr8h8ndPbzPugEbqrImdQ4MdsBU/d/vIlD5pvuT
20mzp8XGR279cv7eBOmaQGLcFHMz4VwMgSaMTDnPkXrQjQvEMp1CfQDhraLkFIrU
0m/4Ok3pdkGLYYWu2hiF3eDPQwiw4bRdFIAKDK1r41KoIk/8fYIG5vYa/t9oxIUx
bHUZuw2Yh01GYid2jwxh4xh4s/BZDY/h9eYjxBiFZvRP3JgnrJGkQvuBkJKby2nK
QXdbQIQHc90jjjskyb5+nah+rH0+4CKnEIgA+JOOEKTz6ic/qlwPrNZlJtEe/A78
t7HmMUKMsNPrvyxOB6uSCZrkmstkseBw0he3KPNas7pbL+ENzWMTjO51DXCCg3rf
jlNMdi+/cBlRkevOblQLwOx6wAFD0cYaK71py/cS5YkiVrgGOts9qBp0Qg8wamQK
K7Z75padlBBZt4UfXuILJhda4EjuLYxC+NogfaPp1704NFL5eiKnTKULvk19SQ2P
tyQW3TNWoWnzkoBtc0dmMd+RZm2q/UyD9OSlR/9/YKcwkI5MwC0exO+XMnL6D4mf
m1oy1GOZbYyLdSuzwKWcqfkOt2VZB3NSKFhsmop1iYvFJxTdjDIvU4Kfk5Pufa64
OnSCZ/B8piv/ErEavpZ9rl8gC+xltG6vIYFYkKddNvti//iqIlztvRaDzHM2Na6U
FkrtQ6nSwG20ZBfi1G4Fr5pDaL+MBJMeplPudMKsno1zyVQMibR5I/ZGIrGPR7v+
lhd4fF79yuxeIjNvLT/UN/m2ZwZbhx6LDbbhXR0WD6m9/jh1ZUHWnbbvchrWkNLL
hqEKuxYGn+qq+15kyCs0G2iADl2ub/aArcnkwzhGoWA4iNg+M2pfuEj9+NXTdYKY
wssJvr5nZLQvtfwhc+HV4VUe2XCapFx0G0/X7+JXwYLnUhlR5XFKf4bpH92PeyWv
GvCc7sMZZGu8/2Cg4bOMFQUHk62Z6sTvWYXwb52JwSSJ+yHvTlO+0jLwQErgE0wJ
vu7aQjo5WeLc77unlHSSy4F7HVJVXkiqW+UjJQKiI/02vS7qtZOTakjQGqFWnd/x
2sjD52MK9MDfOYsPQjEADQuJdsfVEQzut/UUgJP2MkWDsGurRLWSQVPB0FFKu9D9
F5M2rkiF+fv6nIFNDhj5pMaB4R9cCLi/9Jjel5IOVpXiHS0uR0RizbiOiDZINGsb
Y0OLxrTdVpW8zMqZAIjNDqZJ6MEJwLK2BfN8scGnH3xiwoFVuHI44qJ55cyzrIwL
sEhyo4/TBfoY5DHJr2cCq4M1qIFk9UcAb4Whc67Y/IAY99Zc7ioEqCw3Nl167T8J
E/trsO+AjfjjCLzE61wbjoqrKdejU72tB2hVnFaI5iRMjnI3+NHWADFYtX12eWiS
1RhD4mpc6Gc6uE1a6P9u0HkfU7HA/y8gVla5JILybfm2a8uYJIDYtfa+cm0K3WUS
ME7MC/cmxrvjhKdw7Kh2jdX7CRalzsufjXZuefTJcgyGTkgqyuUgYlNhftXiPXa3
nyUtQGXRdq3naZRigw+8b3fvDQQ8IpGWDz5dWmBoZAzZL+kKjm0QbNuQHnKbBIU2
4/A5IbNzD6nPIf0111V79q+IYbgq1roBfA5R/Y/FCG+l3EhjCum8gMPrW9kJsCHf
u0xVkPIgLFfuiRhtHgoyqXp8/PsHl4SOocm0iu3hY53d7j3Yj3qDQQk7MR2d+0d2
11jZqtyolRwtb7lC+9KFCyCxjXoZrCUty7oXcrulvzsnVsqy7/Tq6+4Ow6gqYE95
Hvdit1mbAbFMimJG7Ax5L533qXzMxv0cbiBQhs90K/B83HL2X7Odf3YcDMYrGhM+
DTCjApO8u8ACidOPlPnMjL8puPLkxvOw7qSgDauOJP9dCHnzrb2Mnqo5bCYRLvQS
oEJSBm2R9s/OJf1WRdQ+D/UNK0czR1rLDmfJbPN7NZXzTE8SJFUI3L/9tbqoIhGA
j7sTEh5g3b5eg0UcbkUm9tCmIkGdO02SmWoMicmAnCNOwHOGgMG1V683vMl9MLOw
RJvTSmOvQ7+l/6KnIy3qwRcqOjFLDNVxeo0ef/5ZVk4v1SZXB5IY8ARVxySsNS8m
ByRns5XOp5gkCRc4BNMPM130bbNyJwr+A5+mBo0UMOa6UQqMlvb6B3hdycXiRhMg
xJIONnjLUunUVFpl5gj6gkP75PM6bKkLJ5lIM7W4T2wqEM0vHvKwp3bTJfVlHtIT
uuhlV2dIWLbQb7qYgPkNhskHNTCkTTumkwpWizL5CUgU5HKKE78ni/yFvtuNgjpI
jLR4bWXfnd47mTi0OGJEeGDlaq3yw2kd1tm5yMdgU/5rDAB0ZZ6BhYkrZE9G1M2M
l/15oOSljfZz3GVLi/ihE5mI+ZdXvRVqah0NzSSMbWdiPMd76oNoZlmX64euIzHe
z+40+fluGgilX8kq6akNHtgCzmWv5IQ1ABpWvWGtwzojnPpkvJ7h/PnBPqYzS8Ak
4aGmU+2HVCRa6SYqzju31tjZOqQXlWlVNbYfJSCpdSrR9rUF3NpMjEDLBBVP0sQW
c4V1xowIutQf+gDK+BmD84bnwhPbtQMqURADs5r4BCotfnhjyrFwNdCIQSSpUcJL
N2RN97EdzhDd/PmBrlIcbmojKdmDD7RM2nWbC8YOI+0WHErHKSGFZGPJO0vsd3no
+WGQKhvnIp7GOBDPSy4WydQuUV/KEfGCk6JprdDy3XtO6B+XwZadYn07gn2s/eaM
XH3CZZNf6gb4r25CgomLXdU83GQTkmRlriZ5qOjk3j2McrhvFR1Bjs7MTtOZUU88
DvlgdZ3pfTI3Drbi50kPHMRkRHrU1i3vo6xRFBw2Zpv5lybVrnISNReKYn7OfAe3
az9MWH1njpgJDOCQmDfJQHKJQYM7jgsgKRyN0IpIILrnvS6Lx2o0QY9nndsvRcK8
u5VKaZNx4I7XIxVvCt5+LMnPS/JjDB9Q+sWcguwGV7D1Ws/swdAA1i37AYfbrrVh
4pFyiKfW/AxLn5X21u3iomsI8nN+o8lxvfKI7tWLcjEcuKh/0LCJw2bVgru+SBVb
7tznItxa1g8wsvM5uHDtd6cDsyITjXoTHsqRtFBCAP/BBIsAAe9A3FOwRSlh6nXB
he5K24BWniG8IF9Kcov6FFeTQ2Xrd2c1c8MpNxi8t/01OdZdm7W7796irxqfihLb
LbXSKU8/uJrvN1eTsDF6oKVTAudI2HIEaIghBO1skkRCXZ+fEnNPdsNl8NXtfwHw
fRI3JVrnGFV/MIO2mui8Uu1EfMR5XElgdyglXIUVyvwU4Q0owWnXOslKR+heSVyo
d6DbAufFuK5M7b/ouP4jJPEP6mBVeaSGDkQJrFVt0/S6P/5eciREwTIJtemhUyhx
JqyxOgcxCzOBs+qCwoMNZV0saHX0CIWYRmgxcKk7FmtmaJEmc88EJZTlYNqaX0Bx
CiDyc7v3m5DZLXWkJMmJuFPMhh0fJNA68LZ7C6pnmpGjVsqt0wtPcoNExmEgItt7
KAduYNyO5Dnb22ZjR72QqhF1+ft/3NtPWN5gGuPvAs21yH9+MwY/neP4iHlnV+fd
KCmH3ISICup074q+3X57Ctbu7y/ivh0zD0tFTmj5epKRotXiduAjZt6LwwEuLffj
X4+uSos61CglDgrLd9dePGzxs2FS4NdYUBbVHYhC+SfwqJUO0gy0Gb96npk1JQxH
q+arMAElhhXuhfVRHsNN+IW7rBb153tdHR1b5bO/x90vf8NZCt0H62YgCqzbpj+B
QDWng4cjtzRFvP3XP+KuXGGCctIOshHw7BH7gw8PqTVeEobw4P6WdaseUaZa73Li
Z81x/GdIwYM1AprsbWMwT/o3pJZl0LZ8M195teqDTqOWTTHfi6/AvRQ+/KIa58yg
4otA9J+SthmXnEq6nfv0QX7v5zjRSSODwpVzhWIWPde2yRTE8oykCgbIia5UySMA
avfYdiEezx12zQ6p4cjqtRCPpXMxDVDlYALUmq8HzdrqlG5c8QVWRjiGe9jubOYD
Y9tly+zog9RFfDk+hoNGkxg6jsDukukGyU6TFZBqbzkFpR5m4C/lHMjoGEmilnfv
3OkwlGkPt3Ssct2FmC6Hd8YbnCcufdqZnR6pRRw+5CFRnFwIt2kPmEe6dMS0lZlG
rzhDQe/qafkf4UVym3wYk+txna+ZmuUF9jf7xP54tjKgY/zppzQF9f8VPgkA0TUB
nVnSO+fGi2Y1m/mhjkiz0nP6mRfggQpHhoKsBup1aJrbApHaX6s4aC/ai2hCULIw
WsCJ6yObqXmyDAq3ReRCrzbhgVczkcXJ/iPKYy98uTp3liVa+aW2kJZZekznfdFA
EH82uERehjeFGXKGTRXxeX+t9MglNMYe0KP9afOf/tTggcmapw61fz6CXFrumVoQ
nPZ5MPKfUhKK07dWhwQ7qSMdB+tfFrWmLRilq2FLVdlt57hQTryZ1zruj2QPynHB
GloMJwLpd4wf8nAVQfEB6Q3mxXZUiXJFbxuHMrW+gVuJECWIEjQobQUiMWRg5bTu
mvgOLJAYnu7Veezy3FiwcozrDpuotUfI+9nc44Mlv/8To9iJKsS8krrQ4NBC8nfI
pdpAnFemcy14z58LK9uIx/tX7Cc+o0qHPahxBQiaIlEu9WUTJM/2Ig9vM6JU1fe5
Hflka26Bi/w+J+KCKkEmioqcfBv/QFuXhIgPms6Nc9pxcsUf7ExScQAKgKOWQyEh
uFLeWlKgfUOmGBjolqW2xkHdwXqajFBoLj2T1gl7G8ToL1llccYZEkbyqhurDNCH
WNioCP3xCCxJsGXeuEO3epRlaaLHMu3XVuYd7yUUh2Rsro2z099sbOvLbqJdBFv7
bFsCVwvxENG5NewWD/Kg/JdbYv16fX0BDZlObRfZBy7TGQnW/WFha98VpJsK7cYV
oWZQFKuoR/J4JPA5PfxivKbhuI8HWONUoUzSvRWz22yizLijUeswCZOlBQQwneKK
A8aXD4Ycys/xlqVte2sGe5jSRPWdZsM3kM+6Jambkiu3tvoPijdgpJ90G7VfQcZd
E9Qop/+LUdGJMGgcpenV2PEAqbJeI6pkO7fVoH9qZ5El59MGllJ4Xt0XZL6WXqxN
WLnR4MNJyzk3iuu035vcE1Owae56CwfzcVsAfGmffY4+b5fj9QZuBaFxn8vTGY59
IFA/k3Y3o49HSqpvKOHxkBr/fb6BnYiIQyYWIHCdcEe/6ygufpfexw0zmxu1Arz6
cKxWCDu2S1FNotnpTmkZCbZjTrEp1FzPCvlwJdwqP746rWa6+QjMaf2j5s0eGAur
MOcM9jkjCc8v9kL6D1/RzYTuyO/jyvI9zUMoqEeTqlKljrB5xuoD4ZIXH78l7P42
Gjypwng366ZvfebGWPXkBiKmmC4ujfUivNO+N5j1dk+vvzi8RxoxvqwVxNSOovM3
rIPJ4t20l8omORSkFl8CRm68ieArRmX8C6Iu1PNlX07T9oAPr1/MFtUrTFwy62cJ
7gDpSiPaQ23WzUc54wQr4qQiF2hVVFnMo6FuTwWKCN+JBdQL3u3PEmGs5qnyVcfW
ySWWw5y+zp3iS6VaySSkyDR2VJjnocnRqazNshXUaXhTh+izmIN+KvdxIIirlLw5
2X0yBv/7sV4zj7/ZIOK2fpq3HpVkyE5Xd/ruksbI2ZewvGOpayguDOM1dReHNiMW
kpU21VwNmt0z/vUbjcbsl7mLv6fc3KX8+3sY54C/eXcy5puqb8S7BWlipVM9hpWS
9mMBY8UuQxzNt9klj4dFQBIw0yw30L/U54irhokSEyOoliFHHe1+XNT0a3bJIHe3
KEyYjB1VzVvJWrGF+AgUUeuyAcTqfZdxky+7xpWnf4CjH+A8BcHUE2FFbfSKBGT1
l03M0x5poWkMdBwji86nwDsgPPB+uDPaFSEp2HR/s7dwfOhi+7f1VmMH0oIhVv11
8GScF1grwOxTYTQSKG4xAMF+OCP7o9qgcT9u9sGoeCnXJRzlryawEgThmhLmTq+0
7q5+YUD1LI1ZO8V0ITZ/fMkPHKy1EpcDXmVrXR9wnCXJxOXe5KWFMR3kVcTQaR0H
Apvc+v4tv2jY1J2TT0P5/3FR/DRjTvqBmGxgKs6uaOqcCI1bp16nLqI4VvWlICfz
kUUIULXqHqKbQTr/xtLimZy6IOoALwJs1Imz7ZS+Mv8VQu5etZUPLWhcsY8waSNg
gBdvhcNO+W519N00Y9n/pdOTzArOn5liw36rnm05C4MyETvK2N0/2Sb4+U8LCuK2
4TecJrFXCup3gr3l/KDKOZXsd4HywhTUcTA1cFnuaR/dYX+2xqwpQnfGwa4ugxJq
dhMO1jJ+tUbCpluCrOiOkhcDhn4CNfoJtUO3DUVXZZuJlInh6DopwkP220XLDy8K
oGal4x6EK4dU2PsA7MHS+7OxOgG1tiNW8esTfAHVCMZEaTxv3zAQ8oQ9UXjuTZNp
fBym4rkT6wCd9a4Kf4KjhFZsGrmSrzLNCOD1ajo/2SkC9qWL1nooQFpTPMPPY4SF
U9T9t3XsVKGyqJqoFBjApivYh5Dn3a70/F7GR7JBC71DsrVrNS/SzLeUQDQMqZPY
c9wbB2A8L05qm3zdB2RYev3Nz79o1DH5S28metd+Coe8RS8woSIGrVckR53qaMUL
LDpPV1v62L3beeQxTb9xtdRLM/8s+e7anbjmH6MFVR9eHpFUVWCXe2l/Osqqyjhy
d4w3wLyqsUY/8COgLqjD0CpjIyGibunV+6MNgnQWEzxGuyXUD2ABUmty62ozUHbb
eQDfiwSL3nETV2mar1Pus6NWB9vx6vR0qM9jhyh+fPJBNRxo+68k31SUyNhKD2uW
rYVHJSl6InHcAqFREJ1m5y3b8jV/vvYQrS7GjT4Nv7rmOyWEhC/x/xkky8GWyiMY
TjHkNg7RRHA0fYhyPFQUtRwqwtjWEyJ2w7cYdTfFnOrzHAAGjrj0FH7qOvRjjDgD
GAeGFFCTFG+5SIbuzlsStBTcuBea+3iPkgajhuewiJFGIttc9g4nMZ4k3zffsP1e
jiiCFUqPyzH+c1UIH/jUoo3uySLq8JBZdQUeKIn9Ov4nce8hXf2oIIXOUGMsa7QQ
+IaSEQCr0DvU6VP9vFT/HpRlwEJuyyryWP7q+Z9yLZ8GXGH/r2sPa58rR9QV/NZA
glw34YWSsJaXAjJrkZn0Ajo2j45ChaCu8ZfqyKtB67Zim+vYXhjsH5B5Y1aQu12X
QtzWQzMuTgrlU0xyqYbexAWPfVOnpu0OgEXmKnvzNXhoS8dmsYTQA8Gc+GsZeaPR
V3ap6liNIySI9/fbL792Y4xua3Jh3cfh3NFaebLSBJVjeI3PnSM31/rpRekRk36+
/jsILsNezeTdV7f5h2sjICSs6qLacEMYwLiixd1LJf3SCaC4AGMEUGNOVzVM+BME
RFqIad+joePGakf5sDJyM6PPcs4rozPJjXJKLGBlH09T3o0qSgjqpuDBMbOemgL9
MDQat8EufRAqvTgbUkxbzK1nn9qkYEhWBWpC0AVJR20MtUoF7K9GMALQQ45vMEtD
HgaXfkPYVUH7ihDfwffdL9bSreQVobv75ihSWr4Uw+0DdJ0wK/KwxGPPXzL3q/ow
vVt4auEC80mMRm7dk6vXMGKDMUnDxShq1Hgblvn4KHOxdil6kt+3VF3IRC9AewqF
peX9Ertt9CGP4/e9oG1Ea/G7YN5wTDSc3+l5ksmszT8iAeWWbXUQgq5gJN92EtQQ
vosyLWK91SzFWUWPHSjfEyCcOdJ2viuNmY4vVcTQ8j4wXPiKjK9hk9pL8TI7EkpC
sA3uza+2hukQF2eFjerB+HyBc6tkcKwWwNryRh7bXq5Y8ZI5S46n3AXevUkQ4AA2
OJrv9g0ZrYcQfGD9lebyRmh6WqclM3ihlnxjbsJw9O4F2XwZI8o3rduU6DmE9H6b
BvzwuwM/JQbMiZT1D8y8KYsMY/htJ6ybV3mChX4kWzLLG55wZHtr7VEXSqYfOnea
1m3qdSLY5ykwBwRJ55jVT59pzIvDaD+JIer9LyRghrQs4aQQPkio4I63z+NYhdf0
8slASz4cubDFPVqBydx/IDbja+zKtn3R9CYM8PQ2ERaQsLbYchIU66DpurjRhru0
6u2Xh3wjPbHP3J7IPxMqUbIDibQErIzHpcA3aCfFocJcb/mwnW6rV7Dzb7PjYmm2
pVMST1tcH3z40R/HcMGa5aKrlNuBwvUJbHSVYwckGZHlI9ChkZC9xKmOXnMhNi7p
cWsqiHr0gb4JSq2ZAqY5SUlTdeDekzbm0VM7/nRG6nd7eObwPEO14fsKrrk+smod
Xj3hRvyH2gGugrUMOamQkAol9+EH42npf3Ad1hBPgFr58u7PZpQ2fte4RalcxDyt
ZhFp6f/jvxgvZKKk47YqPmgPIJqH1M9VJjzOk51PfOVf+XH96hstNkL+RoaPzSU4
tvuQblm2lBnEDOmZhEFw6Ba571xfLlj18GD1blIZXoKNv5gIdFnbVKbctZ/rq+ZW
RzD7tPhZ7widfl7pG4voJDbKM4HnYqfQTe5VNJzzLmUi5yys4x3hYztwfLTBVbyG
y5CKk/4QrvsTywBhNxgKm2fo+p587FSdYCpObxB/yaBkklhAiO2yIwqJUGYJM0Q/
bRhkow27eOgIJZvaHAsBlu1dfaaSo89sTL6Ab67EjKS+b8m+b+ciNY/6U/7GUEdr
4LTy8rHtGbAvn7EK0ULZNM2fthS0sA60KCkOjf3xbWf1ORPB85cmM5FKSNTesrNa
s8Uc3/B58s9m9bZIyEuIf10MeYf/Ds0LdGVgCqs2Wo+im/3u4tOu0kdX2HnMZPsz
1LK24wbeUrql3QEtS9UU0b9WBsOLGZ8uGPDa7Fna4nWNc/52fqFQ8M8AujifUiPr
jf2ilE80FlkUSh0EJbDB98Dn4ozght1wPEJMd/QIRtL+wBKfEMMKYBJBdS3iR4CY
44s3xr+FxZ6QwajFHowRudZJeYe8B89Pg1PPGNQwtggkmmUl428pOhQQ1ILWhhf2
2vG78+6FicTKCyKQSOzyMYzsXu1eukiwD3W2OionCqbGd1pyt1K2QeTG1HFk3Rnx
cbJiRB1TfZCKRqCQW8snG+tuTY14eG+ZWHmh2Kao9YCWxkiCycLUeShV6meDWg95
AOa6Bz0/0QhuixmYuvLWro6pdKMFahx+3y7r5bLCU++E4YoE7SArZNf576BmVPJ4
rvUm4JQBjiVYd4Fuqv3NOnra7Mvbq6Rq6/vm2ueoTmPwP5drXRe/Ul6cPMeGuCNb
inKEHjrBZ9oHVWsxn/JHg+XPGeSuous45Bvkm4dAcF8WPuzRCFPqOGS9Fhs+gGkt
THm37215Sgge/nN2LfsTyndQoF7NBdpRogWwPN/lzEx2q87TfAimggYIh1WCCaUQ
HTB6XmXZU0Qx23gXwCEcLtUqF9D7Uf3iOc4h+JrLys9jCZVutoKRi+WntHW0CjUB
jnetzyQOlXI91HNZH6xFisYQcsMJpyBZ2WAC2eBGSuhzRJ7b2m6hcb4UUtLbNT19
ChyPx7+ZV2wKyMHKPJx7OV8RxdnUJyfBunyHEwql9nR0v+OHl7oGQfK2rKAU5VOn
1keo4g02gp3FItOry7kZ+lvFiP0if4gLVP9ZvUBQ4SufF7002AO/i0X5rB+gdAbB
rT/4Vu7/htTCF5m+DdXtdl62yx7N358QvygUd+rBATHecDMEjoTh/mzYVarQ1riL
PNKo0yfV9a7SuMVhXiS4MzsNNGTMyDhjbeWHiH2VWdUAd3LRCdg0LIet5MOJQ4KX
5oiDX2WyV0mlmzGhtTogvdRiZoKz2G01uiBMAFfupaz/VIf/1UtQfUzCCXxvxqt0
furhq5KIk7phGm2ny5WE2HVHlOAvIW/TmXpDXp4SXj6tbSLlR90t0iL6tzz9QLDP
DreF47ozOFBOqdBNpTD6LIbwqLXI6urnxcdrE4HUHdHXZ3wvp7kitq+tFRYTxSWh
u4Q+qgomEC0WwUtJTpOetcBclS1W0gU9oDP6sfdJAKPv/j57oof8z5rfc8Vdx1Op
AYqgebn+dtdN1Q/QqapOdyow8xfUZDy45a3mdCG4ijLBh536t57qW/6wUJup0KyW
Vwd/qgYQQrYQ9FssXBMT/ym3nLOm91VQkyDRecS01EUp4mWj6AI+L0rFwAeD6X1Q
rutyLUV6rzVHNGwD7pvdEIMRmJlEGj6O90oMkf0s+6MCf1Kj1tELE98stITPsBdQ
5aRFtDCNeSkw7SZqM4jU4L0OKVUt2wIKV25G/fqursRTJpEaETBi1wsNPDvoNhMl
FQBeuFuaFxpA5Ps+z4W+GnFK0YejbDtCDSFG5wok0Dt2B9az6o9lbym4xn6Zigbg
YFWMDbZjFiUZow3HegU/4gxpE/tMWSv+obH4b4kdn5bRVlJl5MDGXRasv28rCBYe
VYkKjRhCsq8USJ9F0ZwwbsL6xXUkNapwu4O87MXJhpXh6zOhS4+5CGe6UgFwIi54
qZbOTqDek6GazayQ+JhDYTMpp+EfNrxFpij64NvZjDkKBeKB6z/9UCV+acrnoREi
TUqEoGzqYi0mMQuP0MsbM//m/ELWTben8yux2rmmDNhlM0dgja42x//N2AXl4tej
ja1ntccUcvUGFnK1nmKq1uk3LMZFhZQFyYsmDcfzkNRHa58RtH6hgaWKk62B/KXq
Y+3RQqqxzbwQCi9trQfebGhY+hrhZt6nnFTm6b6oSDzRL5vIuHA6QIzbsZodh4Vy
MDYYmawovjTfQDo6WcXt99hqKadUmCVyaL/omYayQVeNGcqKnHABJ1jq3hcl27pl
8M0RtnkYlNFdmVByfQyuc1KxI64BrYmzI9JBXYjIjIYKIDepAuA2g8V7yq0Dqa/E
99hOrpsYsDTNvGYKPGOOW5dTOIq8ZYyPWaaa+Wdx4E6FWIAwNGdsb6mkcwXk6pLZ
M67z/TLkTojbGHL16jCFYpQBw1HSwwOVxsSEPfK4M2QHlAaf+7SzKs/R2AYkbvcy
45tidQHTxQr80nDYbZPWsdXuOHWK7c3QWrcMi5cWpEyw2RssUv5+14duZGHuwjKi
wII1HeCed5ev92R3W0NGv+BBB/RDGLCPWzDeHlJRp1U2f6x4QgtpOgIll/F7rWoC
kG0JneMUyge2zuhIKlAnIZblF6337sTX6pUX6upXNvJ6FvdjyZphSprOB3uXPAvP
boeXu86nkYVYfPIX7s19xKN7DAXSmXvP/uMcZSuHel6Sajf/YVCy/vFVZutL2fqs
rOZsNFS9Wkghb9hQCRHo9aI9B9gqjUWuofmTgP5oclVcMBH8GgTc9VgiAOLX5S6V
5CBPl6FjZGKlmrrSzh0hhwvih6AX832fV8apE3Oz2HtDPoKrYGx32GZ0dtqGmBnG
On1FzUsg2J4Qno3nwqgocF/fddU57D1Ap1kNs2SYAECjL/CAq5Qny46VeIvuRkI1
B7HU1QT09CZ+D0jma+R5UBzxLuGgwyszvl4ALacHEFDOPOjdVU3/dNrPs0Sb7obH
fl6Dr6g9NSDvMa9UxycsVdgO7fUB3Xp73DLBVlI9v5FBdDXUamXXPMF681F+RcOQ
E+J/VVLUc73uWBqJMxe5NjRQ+ssk/hAez4FJhpckFBHBmVdt3fv3jJJUy6+KPvw/
4rc/uFgLhVNjDBhdgTyxXf3aUKOcgjGkbD9KHMVzhl1ffdkxoAzG50/OwokoO0bG
Xo9KjlcaoDsfzn3xEhHu9n6ZC78ir2ZafRN5LGrUqJKitANXxgdqJKnAIC0+M2W1
GJvpBmYhbxM3xvOVDwA5o5jDqP674+SDOG01AuFWUBjm6cW6Xhf/L5OKh/ysmKBw
81Jn5udciSVhLHa9dV2rrqhtzXFamtmuT6IWQjfPS2ad7FWz/fDkDTK9fhWWfDBG
XcdQxMAGaWQi2JIYbD4lcVKlPFiG4/PJxTjBB+t33UnkGr1LkcxFO+4PiaKjI6pC
jYqOhLAdadPva9vJFbc8VfE3vFv3aVMd/b/7W6kTA9I3R5BJTdECU9+WSZX0BZ1N
Ih4BbI0UfXUD2XRF/NjfA1B6ql4PUbn3y61XWKtLtj4g/ZxBohbUX+n8fTx866hj
Ma3q4IiPLZCZz0FCESrAsyIdA5rplzwmpZwskZ0rNEc45bGsIBMRVOB9pTAMfAte
1CUWsnlr+vXxGiOuHJNm9f2hGb/mgE3SoS1Wi0QiuNtAJQDjeevv9W3iEusRApNx
Ltw0ylQy92RoZNrjOyzvMVdohcmMmSq8HZacYGF1YtNx30Asu+JvjFbTKTP+CMMW
GaiFEnZIRemmOZV12QdVlH6xvfiO3Fe/0gccEjLYmaggfo4Fzri5T17Oh2RzAi98
p2RhA/yyuVN3jQSOI5FH33oLwrWpvr1htq4jcYBqx4iNawevT6QIMhe0J6whNjRo
Hmkx/KHVOfnYDdcAMoFB34x3H+K2txjAtCJKarKJSDquprmCInw/fctlaR76vXQP
JqeDbkW6/XsM3uRBXswVRGcr8mj1JcY+y0cBVjXq/WdY1j2h0WtETg9CeXQyMXb4
nIptiJJoQ7SQrPlDk532eEdksuASKmBy08BxaOiTxydIsBtBItyrAZDbbxAL91eM
WxoycQupPRrC9f/XOCRoIoHVf+v1B7GaR9VW3Dtqxtuj0Lmkyotf9fG43HNEF0A0
aC1U0LH0W3tmBjSXvE4oKszCkeNEsi0V0ecXj9eGxwynunF4jN6gmhN6+TMKKED/
Uy+wc0pjjIFyH+dvNZ1BwAXpe1ijdJPmElJ7/sI3O84cenfpvAMRXSD+08hQIbhG
VcZUgWrQGL3y9Cwz2UhXDBSLGI6F3UeOvAm/S3e3RLzoP2MS4UnAXF+DADpH55gg
GzsVIVVmMPkUZWHZIrTgG0OuQlj8JfE3OV1l1IbrILHAxGRb5d11NrsL5gMm77pk
FOdRAHjfFjdAgrGvmB+bopxMoLuAiHl/nFW/QMw/C+J+mAaO4usnRFI4oOixHWHM
HOH+nm+By2RRtdrEgd6w7+8cmfvJJXwewJy8uRZ57wXwG31xkJ7lee1giaP/cZl9
US/j5asokuAVEfHCpn1UM6TPYzuB90W6B0kZ/KL3Ganx9epP3crHRKRCK3ZWb3VF
AD3ZgEtORpjtSXB3IcFfSJWkayl9VVShB1osvlpCAL3ME+RREYqytzxgXIOiTd0x
5N3hBC+zX0MK+P3J6XLowAtSld9Baku5HQMUBawJoInsmGrg1dnTCFrZI1KJXdsh
EfAjWmYON0lTtv9v/XVndLmqAnAlU0Y/3JMxiZORhJhiry5k7lr9afzycOTm4VyO
jOpjColiUjD7P0GF1ucT7iydLoxRxHaZTTAK9kekNMZNEy1lTikRUvnc2wwZda9x
cBpqPoAhc4BiXpg0qCQ5CZ87TYu+o1coe5m2nrjBanumcL3WhKHaeDDAHxdqNxlE
v7buJlneKpLJgNEoD1gAqsv2z2xvrgoTw5NPi4zvZaiOeouZ3uegnFaIbI+hx2jr
f5PqNRHYh8p4ekJTKH70Yb83PGaeul4VSKlXTSdUIPnMHQemhCXMRXl1Jw+bhaTE
7jt5qG+x9SEByCdjSyHxQS2XHLd/XHZ+Y6FQne9pMZi7w7Bi5RqM734B6OoFufmh
dGCvTjfwqYjabRDIVfDERybnTNTQkz+NG3+8kftYs11dPvIVP4CG0JdWJ/tBoPhl
7/sObTNsxLJ2/K7wjHi+ydqDzoK/9VyS0sGSrkZl47StdUdckhMA561b74JsNX0L
TgMJXzkRNZrWDG767GzE/aQx/SVbz0KS8tPrvQzVqrjMTZwfIKhLWp8EHQ/TfL6q
aaF9BRoHOiLdyIrz7zjJ2SHUJa7Vl6FmNWnOVM1xqLngeeKev26GG3+/Jm7+nwC3
a0Hlj0LDZjeA26Kp/yTDGeV1AK6ne0J4l7JnUoBfGMcLpp3fsb44F+BWZ2DGn6Xg
1fMiAg7CEcET257DyKELojH9kLRCXIOnxThmh/9pH3KOVTJy85+x+1eKpzrweyFC
SbKajLPnkPMaOjXeH6ncGB4f2A+dUB3AmHhoLz3pnvJOHDRg4uQ6V+v9qjlC/PE0
q8M/EMODrQVoUB6pHePUbU+P2jyA2V2d0aX3TIO25908OfJNHLXreZPPzXs0D4CG
5Nue8IFJvmH0y3tjzIWvVFMr7YOBmORysvKm4jE1hgW/YDz9ZATvw183bXX42otN
+G3VhbGyr8Lj87Ra00VHsTDVf9ZoYb6BoEKr90ec0NHt/L5+k/MQsgGuvHuoSauP
TDW0ymacNZQlnkx0X/ytgtmL3o/bJFQR4OkAX82Va218Ds3g/WKl1L3FLik5lTTr
h8kSHsLbetPHllew1ke44BwQuhIHryfTCM5I4auEOCRUEinvguJ7H72F4Szvh3vC
ynD7rdYKYqUhlAvyP2jpwsmpj7dnqZ1Mn/c37DB7/9k5VskETuynsxBGrzo4Acqg
7FcCAzHLdEupvsNghGnSNRnxw85Mnlr4rapYc65zrU2sFHwi6/TriaT3zm7qss8s
SKh6YL71NBx0EGMknD/V6pp9C2e+R7O8MP9MuFaqfJmxrw14W8Sgat7pJr0IJ+Vh
znZ+fDYKw1tt51RRU8R2dERZ7zJ8NHGQYVK7zMmt1JDT2KNSNC/fnVvWE8QKL8Dt
fikUBUjO8VWxRIsjvxLFiLbU9IBGPnEwHe4qCJCf2FbPER+FfYki07l2dFNHWaSn
4mjGvUmAfTObuwfZx1OzNB1DqmCQ3vc7o5fiUukfz6Kk4fS22VNk1+zBD3BfdFiP
TLsW8OaSwtEbNDCR5I/MtcyBl0ZWsbmxFI4n3F6IlTbzpb/q2sBeAZ5aJHFeGIu6
AnFLJfX2BO3rpbrNLLAtszXX6CzhSwMhwxC8qOFK1J1VWaRpAHa2JJfHpyYjklKD
9wDPRtpM6A7k065DIVdtkwKDTotaNckaSFrA8zwNN+Z1tWqRqS4xNhpX/Zub3aGp
G6WvVBSEGMJGABXIhxLMpP6GwXu9jt2u5qIjCftsfNYyPMrJe5dUdQUtqGmqT4BO
EDKyPI/dsvynDrzzDEt8fPzwNzY0DumK6tjfqK+l68rGQ+C7V7Zk5QtZMBEt509F
Jk9kmTstwG3Ogm24DwRiNmYmKuP/QZO1ar7uipquDEpvm4Z4fUFO49xla8HYNSCE
e5/eG8EnxWhMq7T+f23NOwjY+9g+u/quh2MkNSK9/BPjemka7W50U4S8FetEMWyt
Yzbng5Ap4ORLItd69tbqTtvfBL09QQNtyPROysOK149r2Adx1OKbxkKGKaGxqLNL
ZDFAKH0hy1WynCa5ws8ain1J+p/3JTNr+OEfa8D8qgxVOPlGPIHo6Q/M8nhqE3R7
jZ93YbRUj2LHbn+wWcaKZE9w+vYEgIqKAQ8l1WxnhA7xz9NnbVwTKdDikFf2Lg9P
a5aSbIZMWNWT7s+KQN4WS2JBkAGXShMxoYVVOCuEaFFqybQrvXg0Ow7klNpXJNOz
g+HQmB9APEfbAJoPDmpEsSiuqNKibhaIyV2exccVYseYyhGuauPBWvHrPqlh1b0o
8aydeRR5bb8O40CIncE5y7uFyCiTSMDFWTA6/vXw66Ym18FLcAx6VtxzYWaJk6cs
Rf8LSmX35jEb91Rz+qE2gmtbrU/qL/ypWrIBeg6+2fEuiF3IEhvhZxEMO7aO6pGu
dFhyzonFcijSFslsU0pzBUKwNBUBQgi0pUEZKSTRsECf7qh3Ap0XMnvl+FNV9klN
xymY4c2tNsYfsbqch4vbQ7x9gg+KHqBAlH0G0OcxWOGaeNkQXnYTPifv241Fl59J
UPcD78dNNOhAUjdBZExpXIrAbjyN2+xicXBZgG+ykl8SHF8nlNj5L9vAf0hYyzaP
uwxQDD9rVm2rCBeQkyhQv0mBz5qMSrGlNbdlOllxo8XBG60025jgwT+t03Fg9nzD
66xfxoWBznW46Hj9OgnmOcuA1AfLsT+NEL8X35YPL22FKFUUpBosyfqy0oFHE6bO
5cTixKwRqp7d+AgZx+C6RZlt0fqdm6ao600v0hwpx5U792gHGjc9o3/RkxCSl82z
eEPf+vamoaySU5u0xI+Hla+WoZL36WU3Ian6QAiaqRtv4UCpJ3dnXaF3cVgnC4jb
Q87ootHYtx/lVbWfV7M1uFxwSble4kqgPlqBq7OE829NNRiVAbPQyAWOe02Xa4ZI
xy5Q8gSuh4AfXEr7hCY+vnJN4/T4RxdGBdrWt2d+Adfi/UOQ5JX0ZjGx1PUk1ZNA
DiP9o8+U3ZZhyaejX6mqQyEtP190VzJWNBOqiR4jt2ncou7oFNxn6BcsudQFA50W
DbkYAxMhU34TGYgDzr1YLpPA3vIHPMt99Bjq+GL7OmZMbNcqccTPC1DMOOydCe2z
oEsS8DMWEUdl5WlhQdj5ou985SG4K+q/r+Af/9Pyk7amYefR96JYODibGNsEBWKL
O2i5stCbEDmlpXW/G28OlLNfXlT1OA6e7K9Opf2os4g1gkSlRSpGDGauIFCA9KQ9
EFGAmPePqLYeYoD8ZTrLPx5V1YKlbmiBv1YB1zGFuuyFIocqtc37ZMRfYMgV8s3Y
7UphzjDGZ2CzHTYsirPZqmJYMKewUZV6RCy6nAxj5Y1peDEJu/GXh6Mg1yPyHTwZ
HbJsMOxqkJx2mztK72cijkvfYZlgVnF0t/4Ij0Zy6uG1bKFGviQFXlmuW4At1UYS
nhQTfS4HHFYvK62psGDnU0u7BCKZTfB5ngS7WjyA53lM17UwWtJOwJWlpxbeOrMT
A8Ui0vuRoJVxFVxrNGD/1IgeZ8UJBc4+chxQS+EI994hSFBvOvDFKdKVonMbnthV
3A+ImZyXJmmHpd8vXknWdI/FS4SP99chlRP2TgeKI3ebRR1VpEd3lV7Dmj3UldLC
8EvKsGt+Dom3Q9XhJCCJ0RqDQWrwKkat1zeyNVxFUD3WA98kvWFweZ8wstJTOPIp
8Lg7gQHMly1mOcXv3M0pEr3UIVhf+WhYG+GQm84Hdkt9Y84D9sNfAWerAF4Efsct
4DR8MYe7q2fC1+6BC5XWcQxb2mwGZrB1WzFK+6p6tt4GO1sYWDvdbA9W46vBiOgk
ev4uUwwA1+QuPniXBIL6F4GI3VY87fzDvVLb7voQN8ZHBxwTbm+0VUy1sxQH+wcq
YuD4zWusj9evMUrRmTxyKvYhiJjyND2B3ciLtAw7YftU0wl9TIIzeATZkEcMVqSx
fuRwMnzyeCbVOyXxV/KS1+xbqMGsmRixlbIdEjVyXXG8Dg9vLv2aUq3+my9Gos9b
IBwLPs2zlyjqi2JANaKYzXBk+jcDSUcjzLfAsAhVblTGXBT27P+X2siYjUyxlaLX
kq0PPqB+3Ap2D4o4TatT5m6oXTwSmDpgzrgdrDKg7/SnpzxJP1YOPLfCGNmh2XZj
m/x9/RFnVkRUJE6DuG+di3HyyO9Sg9trM2REbHT1WC1xnv/vcQO8yqr9BKaiS0OH
L6Kb/c513Yc64w5I9OKvkuU0yk8+KpK7jkikOYsa9ddx9+2JYhKoJiBMq2SSiepK
Fz2N/syt9xK/QlIJCaqwjOcYoHLXW4dRi5EBvLj1uDgrLi9mFZtC2+eyXbfMwHYR
dBi5vMPBiDx58FSVVUdbv72G2+B27Yx+PJc57u9H2//mngKhTsSaHQWhHkoPE27v
K+KB1obp0OvVvxzXEMCaR+Xkv3FHUkcOe1jHMZGAhcFREotdo/0W3FYyHkyLqzFU
IuOniToC93ks9VzwY2mpoDaUcIk1o8ar/K++KCT9tVX6E/uyu22xGWjT13wGzKM7
YO5P5NdYSuo1xedrOrNlGaIvwCYk2ts6WBpEGz0msXMgKnD0oo3yDpduU7xlkb0L
CgbNjjZ7VFxlmAdvyPLzBanEILR5WR2mFNkWvBZ9a8i+o+obntdmdgXqQzUOS/cJ
7iKKaXBmGFNWSFAH/9uVh+xpIXps5LEycQcLe6H2z5NcpvYUV7T1dJW+ZrHCTdDv
4xFGIwMZck3NGUEYv5lRvuK6ce3CJ3ZevdQpyHKqBelcRKvbAY0LU00S5b8Obhvg
leacV8pgC7ai4ckojDovu+VZ4PAFgh/udk5/Qrc/vXgDhNKXB6vslWi8yAFZmiIz
G6YpUrAzPpx0D6hFZQi4Z9WxJzz4O8rVJRPTescfaBIgx/XW3ONzQPVgzbKpOlp5
60VfkUEwM8xwmpyFFlxeK2wODg5545iDY6BzjJ/8QpxVtacWdB39bQ9oT9U77yxt
YXH5k2Fvtg4NWK63U7RdB4qT9uSgzmEWW6q7CdNMhW7cL00tjmZhN/dO7+ySA8C2
+q0Jdu7Y1E4HPKHCaTdSLEmAdf2eeeD5SNXXh6RT48crXvS7btByq2R/18ephfLM
yEN/BmRs5YJ32TFAumlYnDs8xbhljXA0XZMxNhUQOPESNlM9B6E8p0zccwVqPM2S
daM/qm1qsvuCi2mx31shvAdclUKxscpUFxg0lfEZlnahH4ic51DJ+W7dXVwrUIOK
4IpSUxunmhFqQD4yVhmZqxZUk9aRvYtwTv8W8dP509/hlqD3Lnq2wbC6TkY2y4xb
gUkTIgLfzXg6uy9DukMHS6CO9V/A9rFjbf3vmEvoZ2I0GHV/ZWRkufWXnoSARCrE
FsobMyWi4g7h0tw8klVZzPbSM0YnQ1/VsLHG2V/mN5hbqkiKCdsu048Ta6EOV5po
RboOj6NfFH+53CflAQV1V0gGyvkKHYMeK1Z5tQpWVELveLiRkyXXi4kC2RLJIH7J
nK6iSeMcHdBxP9R36QRm2AJwFshX1qPCpSixxFTz/X/ZfP9knH/bW4/AjE8hQM43
xW6h2YH+LP4hXV+4QOu4pNdQ/5KGepK2kMRuImCyGxq4SzFrF2hDBDLLD0fCdEzZ
3sX3idNrbbU20DlN88ro4w0biNyd2kaX9HAi+R5DfFSCdYnaYMq+hqkiRRh7DgJR
tOis0jyR56B9TnnpH6Y6IaNyXVfaR5lcqnQ4TZNBIXWGeaGwTnILIXtXlDd6h+HO
y/a6rmOKROlfGIZG45Y2fOZiJS9yiHcDFVqY6Hd6GOdTGG+RxhbXKtjSQ5Qe5fiS
/B1QLBZWgLZxqLPq8cDCRIwGsFdiww8YGCO1ux0OAvk2hvWmhGivLDGtThhZNomw
Ti63qx9Jl+9PUihB8+oBvmqG9iwpUNGDA23LRqlIHRf0EdYneiZOsy8Ndx+jEEbS
hJoRTO2LcqP66F12IylYUaafTizZmqSoLvPtnDSGOk72bcSlr5nb8r9xF3jSJkhX
HQKjxAybyTeiNzMUKfcGzq6E1lInbQX1wG+9zfbjI6b1nK3ocEazj1w/7w85EAmr
qL9oW4QIyB1eMuFFL3JG1B+ubI9z0RWx4J588FyHTyWJxlbeyod6NEU4TOhCl4sf
4NkFs3HXQQt0smPoXOmR60A8FJP9GcxriBN/0KLzLrqRKX2Arug/ak40CKk7UB+s
2vkzkdpc0iGIliaBvvfY//Zo7NY31ULMqdzReuCyPQQN6SCcPQUX6S0vXC5UHcCP
cFJI3q74VJ90Zsf96/65ax+GThycjezDdG9iC5J0grc5qUehDbd+CqyA2fMjcVjH
ty3OyZfl5M48JfIlONq36oNsgnxSkk1FU687orZiGOm6LKHqN3405yLagV60MJpv
p2sNUIShIGECaiTSlcqVlZdcNcbp2g9+mZo4fztRast/RYN2H84M03yEzCYtyj+P
q1PIBrAuyk/QaKgKrSFYEfwALMYBIcIBt9AfyuGc0LUkNF3sjtZ0i16iul9uHlyJ
y8r8k0HBAAFVsOg0cfv75KiCH98F/09dEOF8I+VpluEAAAsjmEjgWx9C4j0IZvmP
8G4lhpXPEiDtAGpTVD8Wy+RrUWWisNZ+I8y5GyIgOBRqxi09BGQ6Ht/QypXxl6WL
t5M0E+ESwNj8Q1hiaABCxZiVxFnr4l+XfdYGshjGluK3LDXYR3lGUwPXBYkT3FjR
a88MVtsCbuv4hXV3ux20LSL9U1FrTH/Um63QONz1rblkKahhx7wHg2fTK1kIJkO1
Sv1PBjz9L9XKGhWbEgKgpjpXOVg7y+tox3ieLEhQfjTWCD99dpFreP37zu/UlG4F
yTnf5imJmrSvB/v0Z8CIWTC3GefFn4qlgfgb3HEZ3Muae7M1oVcfyp4HOR2gW74w
ps3KgPCdcJyLaZQx3JsXhw9nUD0ipCCjNwuGzh/Q/gA6CgJU20jqk54BANfdO2V1
GJ/9YY0NYvghaMn4NBI36N8dR6u0XJ8aYnjAtNh7/ffHzq3D/PoERG2dUoz3FekE
wV1939W1pEjG7fbpuJq+ndmHVkIF6EXvRwmltW3XGOrwgfMBS4XHmwXcvGf92jLb
UU4K1Xw/przUtXV9Y3j3xkENkGJhfwfKTP1UA5V0vYmTSq8ogHl+YAyH7Ucu480G
Oor3oBjo5NLsgfm008ySzxTaJPXo+vCaemSdfc+WncYngtv4lv77FnV/3U0ZT07I
dld5sUAJApJ+FWy5viV+/viNXBcRMT+WGreq0vc0yS643sHnFsZ3jYd+elBb1oy9
pJI2KFL86XT2Ko2T4/c9tq/WD5Y42IkJ5Ljjzi3V4eW/cPaT6bEOZahDtV7uQv/a
knBKu9sNNr5I5uYustlKQrrrlMPV8KO4NLnv36S00xbMbPpHZHozHuLNC+7TH0eH
xrFVR80rB/CqCzgaptaGXpv8noV+FEohTnPeyrjdSK6eEvBwYwMtZ5kvDJNTR0CC
kJGzivlpzUaYjaNUEYyrHhwcFvD/85wBrMfC6I7550mx5y1pElqUBWD6bhmOzgMC
m+3Dv/UCChwvM4qy/C09fMuAi2oLuT0pXmvyeU8evUs87wY2LRYW1F+SVGc2rQOG
zBZbuI6gFi4c3XysQp9uNNrJ6cOdRC6QM2+ACENoS9O2lzt6JHt82+bncoZZZ9OE
g492cNzki6a7Ng8rtMGUOsJbK/zJ6WW+OmjbWpSTjd2ehwIkinwToEviq477pJZd
qfpwMvATaeC5fINCPkm8ALRAeaCMnuV9L2qth98k0TQ+fntjLQh+Mith8efpX47R
lXb0Lz1B34TGSuWYhp1AVz2v1Z1DEnw/X57wz29Pkpn8fcALpryZQiLlgk9reoVk
d0zKmMhAB/H8S3xlktj82RPW0Dplyw2sdOp4yDSRwv1BgZDjPNh9U5Psqu0wi0gp
9PxkMRNeaxaLYMwQ8VL++WBGgtZYnRUM4hyhmSqy3nXJuYV2t3s3/J39JotMLjSh
fl4qV/2cgOhEAuqJhqyXZcaI4sOizrWHU6lrHH9PB/MbCiCNRkXnDpK92PMicqpW
PD8lr303/Vu+wY6MOhaDZvo4ZIF8peHaL9Pj9JDaI8PZHyROJ2jUThkwJSg5pWyu
A+2Qw5xPeHcuDf5v+Wc2H5DW1XtYlJLbCsmQr75/N72HqfTHZu8GhQ7Nttueu7on
RwYP5FzAIZGqcF6EErFeY3Ak9G1nX10roc9wTw0uXETgEhW2TW+u0InmSu6dQhVj
+mM4F+xHo0GQAcXzxFZchSqOiJqUGCAVL3oYBgamUEKVaDXJGzLTuJBdkzAUfwGa
BhCfgLQctP6SBKIch1NLfvxDfetK601KHXRSQidDxn3m4FwTfn6H9SrBZHDzuJgK
/OuvaoAWcXtU00KQkiTOa6DRVTYQCIvTtenFePrbmPsqVPsV5XsLLurNsgLBpHTU
xKK7rwwzUbpLKOh2JALj8nJQ0PyYJE02/9e+YUZwxYJC5/9nxtkTUQ2xzYdQ/sJb
aZKkbdnBFECdxJGBwaEAnlZh0bqHdoa9Fwl1h4S9L9F2G6GlAWtsbzPeP+UYXmRY
e/VNogy+bErIyEAeqYodr/UVJkvwRfUoDJJ4enaRXKM+VQUNGC7OBGWzxlhRyrEI
TrqKtOrt5mnwcdd73RrkT6IcC6m1y5ApxjxsAMbltUgOl1u9WTLVoe/lFy7zLwKZ
eu7DVGnZ4rQQilvQPdQQxzXpV3bKL+xgGy3EZdsJcRZMBGoII4+yzd+K5YksdxyC
0nHBQ3wRyG9XkQ+NZJB2Qfz/R2RX+KOVuQNPH+2yD81XKm6D7c5GZ0k99VWFJ4SC
OOf46jj/F1q+bl7zDOcRE570ZAl4mZ/efNUplJY0I7CXjtUEIeHEl7cA3YE7d5El
vJnmiDUm3qDNU+2PluTip93odKSxFbf2B3WtFicL2rJQ4VrYaxl/Ld93c2mrUvyF
J4U3SbpxSFaQHJ0tLkNRZJbxpsJ4etAjJdoz+vuL77SsMMoAT1Awc4p1XDpfNYAw
dDWA7UNdJg84PaDXwNoZp/X9RvNGYv9+2Gt1fdjy1YMEOpfW6KToEqWmG46YDJl2
EytBMGBRU/1X4MQnSxidnRi7HYy3asz/Wn9MpZ4nkWvuUGdG3c6fTKQ5W6MsXGDP
jCSAR+JJ2qcUOLFvY5LIYVD62UzR0vlkaJbUL7wTAvDeqUfMZ7BtnxtpXAZmlH/T
mIEordCbczwYjxpKUMJZgFkC4rTx6+lyT1KLsXtbiq6316Cq2R9zvKfio4DW+O8E
vAPvUvIzpu7daYNffgGjvfS4shlfl1dRhHOI3T5/Mpv51DWDDsoII4rFNAi4Ykc6
VdoiIoauF/h1bTMiAN6tPwx4qWUhaIpgXcnTg8LGtOLVLp5Y+9Tm0Hpl2xUD/kAr
AGwUsrurPcxg6G2uzZ4KDIwptw5jUEtzoBfM2VhbKlp2HaASMVcpQOP8YxCsj3Kk
nwKKVRZvTzOX3Nt65cU+XsgvsxGuRqzeUUua2gaGLX8iSvhewPZD2Wco0pgIcKfe
GIi6JEsSAIeDsRqahUUvylcMvkxp/G1rnKp6Z3X50elXsqAw6q+mSi3nFvNpfJH5
gacBp3hhXN3ttXCGU7xC2A6DpAsG1Dp1B5Z7UOQfWbqLIxvo1+AkIoGj6XoAGoRz
5+i3w3f3eN/Xvslo/pA++JC5yEfrf9o8VSnZDgBHdJu7svq/A7KIc4m8fbVNtgFL
4mGzgP/sRj3IVwLLtfwe664lGv1UvyuFbFu4C14P+NFHx4fSQoY6wpKVOfL1S+Dg
M6AEP0xqjoIXgu1ArMuUABF6l+IHJrghNZw0Rnx6w7JJvdtkeVwbugJsO9jEQB/e
UCnH4w1b059nHp49CnGD1fpgUxBD8igHHk6KHSarjkrgTFwioNUAYS32k4rD1SpR
iy0zo9RynWHo5yi2G7VnkT6UJq08R34RNBdDnGh+JOh9RchN1aEIA+473UohSYVE
1vl+0Xpkh/wRBwGXjeqyOja6hVY8DXrmAaIx2lajdNNr6IEU6fcZmafRvtAxZ7DO
hpmqk31b2maEB+MkmfBbqVbzjiLZnI32EPwG0OQ4gst5laHcoivWeiAh2fjWLpG4
YgR/VtzPQ5zFqmHS9GRTpzV/aufI3NhZ/X0oKDCFFa3P1QceIvuLFoVoCaY9D3/f
euEZ+MDkcyLO9IaDrVePkdMfcdvJ2Gesux7Gu+iRjd5sHkhmySCojUkj9kkAg8Tr
VxP+rI/1HoeGE1KBFN3b8EHKWll5aCqctt9OfeKrV0VQRixr4GoxKB+h5nVpdrHF
oVfT+4cYySfxHQxg0qIVlMEDzjBDvgsIAnmeH7ZHJF2l04Wxh/iBVOfxDg3wvG39
G3qdUimFe9n34FeAayMzwycUWkjw+LBeVhj0cYHcisW1Qy/i8TMlJK9gO881RmrN
eQ5l2x3ux9l58GKXSZj2X2JZIP9K3jKFzrav/LSX14C6bhBaO9FFCg1RVBtPTgt9
dXfg9vqqpVunBSlutTIGi8Qk4n0xXAM26qqYmXYjxAfZZyIepHuRqYdvjdF8v3LN
vnFLpe9mWQZLSSqslVo1U8ODy2PPDb4svfOU5ZbLGFLVTgMos/tPz9iFUZQ0MDSh
1zcaP6874FfqtGNuBx/mH9QQ3wpgo8hn7PyRATYfHyR0JD5aDya7iqMT0Y6lclG9
+XtG94SZbfgSWhMt/fD0IRyCx5jiZKf7TbNClzRm8dgjxWTYdBE17c4GJI7y91c3
bJTcrEGl0vH0K2stiy+VpYrKmaanMF6KFfF7R7iBa067uGyTEcGWFsErVEsxwRjQ
OU9x3+A5vUlL7iFVUWXImSW5TLabzEj2r4p/YRMejDwOyZpfHeNFqAu/OaxK8W+X
ZI/G0ozTeSvrRd0KE1xQ+0iLvkQii7I6ULiueRv5z/a+2X4JLT2RK+cxiUy5cOJ+
oN+GU5+XvaC891KKCCF9b3n14ZIhzs13SPLIYOg5S2cxeRXcnIc62Pu/XcwqwUs6
1dOp7pXE5xc8pPpJRGz3owfGXv0osBLkq4Wr1WwKREV97XC7W0Xp8C6dQ0Z2dPQ4
kIl6ABnws9xAq6Rxfdrwbn6xXFTzDgB6RqiH0OIw46yUyC1VJODCW9PsrAZ5+o+l
TUeSfRTvvaBORG8sgr2MD7i0yZvrjg2jNgHZS1KXHVxY5O3CN3DgEnAqgVGsnXkK
zkWlGvuFxC/8yJ30paLbKmxi+2oEvinA+hQG7u3PF1NxsMjozQURssjCFsBxTJwp
5hMXtRrMf9+zYKkvqEn90mpUEG7uXagzuFMvmdn1PGo/Ak72RCBBF0DH3erPGrC2
NR2xIi5735AyXj/ay1quK6FZ5Uu+g8u6aGqu7159Qjsq5D++Tn0StGIQmY+3/GAG
hheBCfiRNp558Md8mgT7YBQR4yOQfsAR30JbfN8ghC/PXSStTqcmjdFZjy3VFHPc
8i75vhMHo6vPc1YM0J0XPIDrBa4OCZn/QKoDiaENQyymIiJhJhSadn6rWQ+z34QT
ZloMcTAM7R0kV//wdwxUioQeq5uBsAPVg/JdGWcVjO97NNgDJQ+0alnvCPFzf4kd
50PY+XPsSUSD5fdxAn8K0UF7Avtj8E4CBPYxsJ/nN0wSK6fURpL0PdzJRDVuHq07
ETgMsV4D3dHkRhlcHiNNM4TWYr3QZQsy99uaEdOjfXP4LSZBinPc9+JwUDbHs12z
nCQRsbMk+eLmCS3D5agUoUlde+FxVP/1KX61JfEoNv9rpks+MYIeoaWX2fO0r892
6PONzdNJEd9fKZicRlZmDrdgsqtyQ7go3nTr64GsbeW3ICFRPlDOVcF1xPA0m6xd
Fw9VVaWOvToAqlXXbN6o2Q6a+z0KAXc7RwVSk6ArP9TNPstXnlqB2TUzUaEtVfHx
Cmr67YeyhX6xLTxloTELDmw08LDBnSVZz5THBceT4DqrTre3Uzk6ycZAiqayhDaG
ebQ6vchSw2+h0WPF22P3iIQeBnsP6NoVokXSxUAI2q80eIGztRVj/gWAQV9KmqCM
hbdf7Ppz+IZcSyr5SgVqjDt6bCC54ec1ys9jA5GZ4erUAtrydYmQ1g2GO2fPHxHz
dQRbsHPf1uFxXk/8zDwCb2gaylD0zy2aWYU290UteFxD3E9zYsFci1Sf1cfAzeMF
NCQ+lioTfYpqDt08S0uloG05J04AVNoFsVgcNSqr0m3tYlH/hSj/xSDSJymvfomL
a2LaI/uwJpU0bidydKrQjkQZuGlJB0HUBQq7cZSuO4SbgKfxNvmpYD+1WK2LXqG2
S8mAB1O/1ZB8Axi37pmdh+5gpgL/llaUEgdNRfUfs68xgCObH6rFvqM6n6fFXbfy
WTXbyeVs/aRwzk9K2LLGW7JoHzsFSKUuxXL/vVGYSV981zR05IFBi8T7jLIo84+x
qQXEmEFgoPuw03/cXyshXshsEXl3vuhA02a0pfekwH2QkMxpHbf/ytB274dGwxvq
HHSVW+PooQFTdRub8aNsM+mKiOUA0bbcWySzwYp8vWOLO7lldexYI8vkKkHErOSr
hs2bjKN3IKLyWeRGWA5k89yAJR+PupLNY8YakAqCwSi/yJiAycJZJl1uVy+Te2KY
KMX52X4Wz504HYZck3GLtSUhIyd9+3s7JJTNOnle2uZpXNANb8zBltwhcP5Tlqxk
3JCmInTDhwzRniRx5BHJkeoaXnt3Bew+iNbMce/jeUrkNm5Jjtxry11CKr7ccDHH
fadtMwYX6FPn10txhRuG8DyR+82do+JAxV+55pa6jfmNcX7h4alAwBrft9eExNso
9wHTo2HUdz8RTnGXyMvlpOG6IKPe18II2H7qT0XMPOFYAzd5qnF60EwnVB8sqJF+
e0TuKpmqysoRn4AGhdF9Dsi1VTQlk4NpScTtgt+G5PQE4tPh0beBLpVADE6zsa2d
b2oNBD8d8mmKYRE5cWKyXUXNHLeGssf9+VAD5BLYo3ZE3j6mr0uCMyZdOe7O+K32
LNETNQk1xPKAbVvvBmAcoOgNXD5DNGrgdKRpi4zgiTqF8V60N1ET0cylO2kKKXQu
OyQkl/9CJ/MlA0W82E4xeJQSaiwY0J4xkZ3yQ85gzmRSRuuFgLygaz0dyjB7lbM/
hQx9bFkgs24zMsAmxZc8FteVdGQ2YYeti06wFOqeMCP6MYFvVuNbrX7jmEwuFjmI
WD4s/r0mkU+skt1jxdoZzsOluYU9q51PL3OOaojBeB6atAMJo9b0xz73B7U5v4gD
lLIIaRo9CVVETxsrnFeRg5roLOR8LuHJBh2UzDGh/wI0GY0sLLoMpVfQD7v4Hyj+
NTo1tXrWPhrT394BVJk7HwWlW9DXDutAR5aBXefIHSSkrNackbfGEZ174b9e18rb
yX+TBjzJ97PJxA0nb8mgk1oYG36dPP6dR9oOjMPJ6Zrb12qV96wOScts9rctkKxd
ksL5SIpy/4uB0aEE5WFRSWFuRRdr2XyGFLgHemPTFSia5aJ16+zcl+XO/dV3SYbE
0Yu5QSGpzaUc7ZguZC3l8/PDWTe4c+ns47yN9SI5zlg5oS4cBaaMsZrFZJdAXy+D
gsJiXixeliyqsIXurAmTk5lmd9pvfz0gHu4MofMMk9JN71bVkIilZ/mR8rTTneCZ
C80vc5U3pp36p+EvAzQBkkuiOzgJYGfKKr8iVaHrbhUoPyRZEdYHHw/jy5zpoDMo
nczo7VF8nXB0lvuEpcTSN3BczmJRay6Km+yIG/oZE88TvhiNi5esMzJyKd8lsNak
P/a/YM8tIdH5dDcGw3qqKKjNqYwMW4dCLbYZIi/xHtqv1Em4xbTGuysSF6gVsAVK
e8Jvz3ha21FukdpGrIxtGmRICFKJ6f8ZuQ4kTNZBkkxo00dV3zWhdjD4o+GNepV8
8tzzdY5b3W5Ch/FgSNRlUiiZbGsHMJFeQbVZUQhX7d0E3wCNnEzsemrY2yHeAsln
h+LRhXYxN1dWKVb3w3O1DmMyYsp3vtH07xnK6x8yOnp0NJkuKsfIQtyAZuTH0WJr
rv1LWBORwARtWfH6Tz51DWhThqulkF9h0C0LrI0Tj+JBOethYSHvcsy7/ahrn6/s
3shIcvD0UcUtL/52ngYYqSz0TQNdc3a4s07Nvj6pvvi16ruVd1t133zDmt7I/Y+W
7Pa1qMOwdajpN2pgBhUCwEz63XNaevGM13PcWEhisR/ZGloeJBBFlm/uqk0FHgJ5
ph59TRU4hG5PB5/yl38/RFFnyc0+LF6vS1o5Jmzd9m3QVVKkvTcGGW57nDH9TARJ
yL6EKQjWjd5xjNu3OnS9+FRIkha3tJhmUYILig0dIGtIymxUBh/MVO94Tj3MWK02
X/Vdy5/GZiNjSyppEk4YrmeCWp9/kizXYLO/9BUN3OIFqd+9Y64eipdBZ7UX6kEa
fEE0sAw1Aa/XxgPNCw8Qmm/xSecb/MQ6nFwGt/oyi66+47RbP1+BxWvmALF3b5Il
lc06gHR8OSdgEsIgoGQHyiQdGQCpjqbnb4n5/6dm5I/Pr38L2n3aXDYC0WD3a65G
QpihJCT3F2OrjSgdiu6okub+nNPHavlC/ixXDq6PkEPkbwki+hOyX25QhzMHKzNd
c7jq79VOwmNIom9uiZclSQ45MeLCSoVI7+A/gZbl7FTdT5HKs23n96q24GlEIen2
MDVSAEuwKOkvmDm0JtP4D1yFvBFB8TYGUVjTt1WuBn+gVXBTH1XI9rnpZzYm9EEh
KvR3Kbwht8IXVR/aWE9xMmZzmK8XT5/IH3pQWogHpWk4oLmoxTtjQcIxawK0nGZ4
Ye4aAl9UZ8nhCXHScLgMLMo4GZmlIL+uRFge+kXBgegiSr2J0H8IhhS78Jh5jZBE
l+DpQy+ACmORTz2uQR3totF5ZU9WnuThBeCUHyyV3YoHFutNx8J7j69FvnZbB+R9
qTjq/Ien4wb7nx6NmUddJbAQlVAjL1J86niq78KK9wJ8UBV9QmBQXfipLL2fui1v
FYKl2PaHGri2g8fMKveTd5o3rLSD7j65KFpOQtI1YNmBK7zqeo3uZbnnkyNIX/Vv
k+D3mMwbvQOdkYztrFX1b7LnTDD071F7He5AryKlXVNe7tPourV8FI0IczhiCysk
svHZONyo+poWuUpEKOa5ZxF8MF1Z1HATuoF47oAPB3cmSesXB7ILZ/6nR1oX8ILG
2wFtcn75DckrCZUWkOGHRfayCLkS+rkiRv6UevfejiwUhsQ63xEgikJNG58Lq1Wr
iNQ0cO4kCjc9ZsPyhaTyUjhiU2nj2cOmOJUCxNY3HH50CAMG/D6my1QpYcZWTwix
hcluADNLurr3lOnk0U+XcCbC29l2jYw9+j8wY/KH8GaQ3IpsnRxfGRYYiqajyg6U
axQXm9sPHgKvfq+p/TNcUpuoJmG91T0RYAchYOjhEAvtRlQF8e4OTFTVkmD/wxnt
/fX8wbHIpwTzVpIQnXgoUyyaqRj8RuqzSXPNjWhSzhbiG2Ab9r6xHgQH3iVnR7zK
QoEQgP4mMLR3Ej73rUHCJ1Sq06wQyqimiBJoeE15pWnM0adtCz4HwtVKLvY8vGS9
NyxJ2FbtTDaXrGoyxHWKF6e6+fDt3bfa/Nb1YFiLbiX9PEHJH8P9TyE9qoDHamLn
2PPgwYQ2CEMYCRm8ctkZpYYOf3SaS4EglZsEyzsHUx6RWc+ytgWlmHTa8r90Gulp
Ook8tyoLmoTL5YJ/rGUVIV2qOsbp/PY1anu3SCoo9uHW2a/3odSkfiHgFZt9KKX/
nS4QLvWG70oU0jLs28io5tZuAOd3D9sk/2LlxIYd1VXfypyl2vKfa0e4lyl3N9sW
EilEze5NizayskPMyaSmUNW7fruxy9cYScyNuJAtw4f6x9hSymQNf5SBrd/v59T1
tv/05dUsab0hM2Kw/FKGoIY1Dj6rHqsuxjRrP/o0LmtV9mRQGaT6+9QjpE7iUAZg
KQ5kZSxweyz3FqaWC2sBoESG9o5NWrCno3RdIfhBbj7IcAENtagH6C3Thzd3Vkcg
BJ4RzC8E1j91ay0oBFEYFI/GoUvcrO2Mrt3KLtfEcBbEXxYPQpjtVqih+dKbg79Y
N2JuHOsVI7xnYDuL9pSfBlEf90to3CY620NX+jCkQbgyXNjpdhup3YYrllZUcZtt
IrlwRZz7EvvMUYORu1i3AXUipjYGUTj17GwLWpyIlso+Iie4BAsQYYfC62Xf9ZPF
jPJGXHToPeyVqlkSkx7hUfPcOOvbNGSl3Ui4VYxYDVbiY5ffKkfMLDWejA9a6yF6
Ah8OthdQ7kFj/q84CXqsspRnKOWwwEkFZZ8+IETtYLyaM+4N3s3bGUjl6jmkFRaq
bPrRnQcBBb1+9rELSly7pDnvj9euEMRjeQwAT1R7AhRcWHIUf43UFJy0rXNze029
fLkBmXS6YS0GjQ05emRWL7cnQqveJwOatQ+p3rzq7t/mt7pb8LxjCfQwG1FWB15z
omazoBk1m+bnCEvJLH+ifPpx3E2yH7uXjpOV0qpmmfAmEf3hEybn6QS4WhhadwNr
NZ3hn/hTbvopOGWbfsbW2cD1yWgPfOZSWUSpDCuYKBWtYH67roWfAqdPehEYJGNU
imZbYufXMG1xAVDBxuKt92ySkM64vw7D87L0oEKi8o+srqAtzsFQQ0bYEawUJcUz
2dIGuU1Mehfi5vBzK0iQgxdxiNj7dzI5Bnf0sBbHNrtl40QsSp3qDSq7wVUGUH8x
BDbX+Dc/KuNFL0UtSiHAzaTIlsTUPJVbfF6VI3RG7rkfXAmo41EjdbGhSl+T665I
+5oHRoqVVINBlaLDLLZH2i3Ooyql5CTEpsJRTFjWJk+1urxBAUsKCvhjzgRkxgv0
/MeFOvmKvkLptbd1Tej1/X6dGSpzW8nuBguUhBtAsyqQjjzyUzmKdFEuh4PoAJuj
DyjMi3LDCa2MCYsJuI0ZB+QT45aKHQGjWiAGo7kX9k4/AXDLA6T4C35laoTzveR6
QElYfmmH6X3cC186aRBMBqE+8Nz8r93i8aAxzJo+/OPXGaRC7dotfeXxMaJKyJ9e
msbxvpmm6d30vGLy++SCVxr/jK948ujVstLifHHUd1+76mAgum04y3MA4dzN0ePy
JWNcq52R2+Ro1yUQKEUwCNZ4HxvmWQbIUFKyWQC4kVGtGWWJyDvvpOojQT/nokFb
FrqGRh29rTppqH41P34cMr1vItRZ5MNzURTA0UYigVaHayMphK9BoqA61nJfwJQp
/quyknzAQa2mC9vmbRepnSwTXxWnVLPLG9B1A9avLffNrHjzlMLpRTjcokJpwABb
8sJIkQViOxSUPvcAvXwFKCUiOfwJJF9UB11YoSZWmsVQaM41+5XHfVk0Nj9uXqNS
piaLmheAKdZHX3RK8Kx25AYPP6tLVEMXXmBGMPY0nCclcXeZ8b5g3jhoq//zjvuX
Rd5Y/HFXRCZEPJiRJAa2qugK+i0EkbUCfRTL19mXFYufJLsokgZAY+Fz6pnRtR4U
izsvfBq8U/PsXdobQ03cn5V+gC2XT+kHIyh9wPMZpvdGvp58OcVif3+fBs2hQE9G
+Nd0SYGJnvkOuZVmRY6A513xZSgu1ELnEDsQAobKcK4QQPP2GZ7Knot7A4+c81lH
3Au528273MkLaIkD74HS+dbHaEInIWmg/+VHhXkj37ZcZeynO28BEtwkbJhRvloD
fRE0A3pC2DV28Xd3xosNRNuMyj75+QBEf2mKTpfl5wB9tcVh5kyK9gUWutn3QqWU
ESXlbwvFyQOR7g7ZdbgGyu2B7rrSaXh2x3pMJ45+nUSMuWAdsSmB5UOeAOmcNDRG
OAM/dEVqlKhwNfaIJRUSYaROdKaMJDgpBjgS9TK4gMkPEadzP961rBiBEzkXQYrD
8HqZallcXGut1WSHoOKLUlblxrl3+2o/eXtQm/YTlXrCGV0Mo4g70fXD16mK2THr
8yNs13VQqpPHOQq8z9cykibc1OoFPK3Ezn6f6DazaaugaIf+II4nmwcIzPAM+vh9
5Ekm7tDPjPWewe2gDyFSNtKTs0hcclhcGWVBEdSOLWQxg7YWhCH54N0yQAi3tDWJ
RvjBaEWpezgkuwWTqXhHPLtjQc0ukDXebVbp2oNozATCOBwR9TBeQIVOzNKlSptG
HUIkjwhfD3liH/IzqUUfFcCuNzcowKR0Vu/ihWPDzCW2bxkfpiSSbRgsa+gwDZq1
333r/f8CZb7JhyQFEHrf8rlRrX1x+jnQJiaax/HFWvbOj44oJ9jIsMtlmJ83HrYX
4uEBsSXMu+Wl2mNcAnuni9RPjKo80J5k03A7w7yFuHtKk8eOlI+u921eiT5+oqMc
vjWLuBojQhvb/eFp8KAerDt7EUPEeTv9CpT3EaPEjK0kmi7S7dMg6h9LA7E8GFh6
JJm1Ii3JT88WYCB19PozzFHTlQVUPeU9uXvUYnT7iW659nO7nwA4dlZ/1os99F5O
2bM8qd6EhACB2CRYmiYq8uusp9pWtyvwR2UXVyUNJvTH+mefjMl38NZgM7uQj05S
/7uTtUZILdS2ZUWRvIxhf3XiT88Px19XC3glXS8YPH6izzUynM3JP+c22+VBeNM5
N6PN3jiEvMttQBAoj86mv1pdDNNrS9wPT/s5Q/NaGZnT708LzNT3hO8BEvpYZzzS
P3xiI4/gVKxgzn1tTOSAZ87Ts4UU230txy0wVgCMsCSsS2SOrLkbNArzSnsrpFwA
m+u5mL40JK8a4znURl7My6j9sDSUnlfFulkHT2AHSCDUgoN9iaiNpRsgNwq4aHPO
xsEhhu88M7tbe3grYmIE4XJzYXL2Fo1IkzK3J/q3CbhgPE2kSW97Z1sMMWgiBfLN
SZ/ApwtbRFIDD328Z8bk8u/u21L7HB953j8iIQ3FNCGvFX7sDS2BwLjyxkalQfut
H8/jGPcd22KJIuFvPjKXtYWWM3HrC1F9tLZ4QhdaajGhxnQfhE7GBsPNMd9eWLU/
+zTJrWRTDbq+QroFHVxFQWVOTy/8eKTEN+TFkiEmNWF7i6uyPQ3tTBkwsrfsSGBV
rEU64FtKoFeZSf4cj3K+eCJxkOFfkCTJyXaAG2i75jdRtL59Bc377z0fC57RMYts
IsWFvmfr6Ia90zz0CF5hQjzOasuQZoLo0x/qag0xJV4WU5ak2gun96HYhkY5WB7W
QTSPDYvdYIIMX9xhg9G2YqmnuUewE0LvfqF2irBXH142wKrYdxC4qOoQkEfvXTPf
OIEfiAItzh9VbBlwRX0rOJf5KmN4Zcnssjwt3dwZsHmBWLexDtRpyE1iPWdFCRmQ
571ekFzTitwzkoT7nxcYyg9MS6tkrWCrOhPoYK7iYL+9REaAR0AR/u4Ihnzk2DD7
1SDBmilUc9wNJt1txTxkBLdt5GP9kRXmufa6G0r3Y1wDUKA0A5arTtoLJGqrCjQi
tBoW46tF0DZxrxOlg5wOdEf54on795Bq3uESUgki+/qIIz/CjtsW+/7dXx8m05PB
f1Caypjv8uJLk+R14doIGr0AraJ+nM2221p/IwBV/5Vkh00ceciDaYFVcXrdwRbB
w17Tc8l619gG5tS8Zl4RBX/aZCltyKmkRefB1LjCNbyW3U2gDs6E2TDW799GPFLn
2PZtbRT2rJyKXJPWJNse7IMMGp2Md6t+jimhytGTdKOzTmkzHipF5cTCpFcATDe/
tXOmWrZolWCsj0h8JrFUGKk8mE5oxONFN8m9SYwUxeuET+wz02bSj+91YLM/BFAT
MTuhCmnYN2EfNKhiT1g2Z0hAjMwZKACqDD6wR1Cuy+utnuKWnmLhdm92L5qUjXRF
uTVvx3bmrhwn2DoReGg0fyeQa6xLeX35roY0ok5Gi8m7o2yRGRlnDiN9ouRlz6G9
VJ3B8kf5Mg+u/UQanMmjH5akX+UYoBhJAYqboWApqi5bWtsSJ17oxigs0pnFqD8W
Ze+htZ4JBrb0TINCvt2eW+TQwvn7ugBLShrpR+RwOUteaBmZ0q15N4aPyvYskQbV
pmxDiHNV7h05afo0E/ktFVvF/c9wkam1gK4TAYfX3hsOxeSxGvkFH0BeT6ZVSLon
5nWypAAzPBGM08jj+rw+SRgenb5JHq9vaRx6bjo1pk/LzUE5RtsM/JnMWP6XApA3
vUDo4FnXJg4V/v0u7cknQdapOMVPJcJ50m4w1UnF6nVi3ZzA7da+fHQw0L4D21ok
ZLjKCrgEl8Br3H5JsvzhGCNHHa/uyMGZTilXUYa8XIqhWKZQWT5kq66YYu2pw2+T
ForqUHZN9ksY+zysB9OsCFEuvWqXXDr92TrlxGbVd5Cb721EMsVMwF9Ztpnervrz
IWQqqB2Klquql7ryKX4n40Exgo4dzYmAuvE0nhQtRa5Srhncgu4x/RXA9uU4UpH7
Bm5+tj6hLnWXXyqP9BS+aZwjK0R0fpIJB4K2Bxba/Y4wHX8wAA5WGuYoFuhJz+yB
SQ4XGYgsTtd3fKrQtRa6k4VYrqM8NjuHtUG3qVrIYTW0Chw4ojmY5jMeU/7fjURu
l2J5NrvhJGI5cESbU4lPdvNiQISM7efyDbssk1PfPWG/wDi9E8YswQr87EoGJB+t
BuU3sqBVKL4CJgniK7my1rJN7+DerUbnjVxSAfvFoM2dnHqR5jYV0PerAEBBWkw6
yHAKmArOXSJ8rMDHJqVLA67Q4W6sw+URQTqRKv/D6WGd7+oq062HghT2GK4ukBPq
AWJZlnXS4yjKPCwnVZJpYaA9xmWQzpWkFFxnsCEgSFN1XQG82GmRYhf8mEOeaRTI
qfDa5E9Zs1eSU5GTCbLVTb5xiQwKMHyEJrh3YNhfI+ojU/EFlqgItY3ux4xEjI95
VJbNq87Xip3k+hozGvndiS11yzpxQTkpxCvRDfMSY3vpnLNiZAZBFFNkGiRWO0Wm
dPnIUttnA8MIDA2H0toSOggJqhSYpgxdCBwF/azXLj6BujYSf8YT5Ahsx0H35lsk
jekeMSn7++7PlqARK4sXC9hbDIOBEgsgwFMq2Mq2A8oVjOVInu7r2XmXLbqmTUqk
jpSkYnujz6dfDqVuY37QT94aGvnhS+aG1k70x4JhCvmtRZ/bd0urgvnHYgTqSqGd
jFsvl/h7yNEjRbNg+jLmxXVVIJ9HJsSoKAfpvg9POkDxRBjBLxGyLTxn6GMfR8e1
hZUJfrhRhQ5m4Bvun/qqznIEgBwtkTXu3nqdm5SrP2iApkDFBDnxCf01h3SUVh2B
sR0kimjikf+C6naaLeGPawexWUlpp+dNS9xqk80Zs3VMh8aj9TMcojNWIfT4aAOV
ipjZxqxabLlYUkZvBLD4NnUqB67r/5Se4tY1NM3Ejy8RXFhnTLoE6py8SvMWsEL7
P+M0ZdfIrYUtuKnXRs0TzlIqWT5/MDFCPRJjkgypOYSVBsjJyPWjIgXj76xeeAuI
wD31gVlk6KamB4D5Rswc9eCwxoiIbINjCOkGOTg8y//T0X9ovRUSQKToEg9QNLQq
/AASqPIGnHT3Ky0Yrx5aeuBri8sLuXcECrmdblt0f1gy4kZICI4I37N5V6BJQL27
wHzulAnvyed5FDzWQ+sl69FJvPXRZXJ45lvmKQh/+otFuiiRvxSdrMAUcXKig5du
Qe34deSYEkTzCnJNCan+iTYT3uX6GRFHT2KYmqjTbqg260j+8KMqu1M/Jeb2a8By
vR5byW85rCraUG12EtVT3ZFMcl2NPo6WXZ0xo1AeiLmbWtM2Sk4YXd5E7hHv/Xta
7fdpTzGVuUe8oYXaacNOeMM754FyVKCLh5XRmOYDJavV/Ssfzaw0jrtDoym4tJ4x
TXHEfVdvzy2FOAHROCxazqBvgkwxakcR7/I1VwY65L3waARfQ92j5DMFixhAt8cY
Hr3x7D6UcxUFGE1ZKdlgg3bNm1h4ZYVdT5tA75/cFnms4awNv+DkS+EreEcVI7Dn
eNHqyJUHbLVjqglsIFKgO2pAMie85tysLTgoY8H2tZBRhcevxuCUMniXdkXBTDhd
YNTHn+UFch/posjNIlbY25HO8IDhA8PH7lrXXzXp5iafyc1MU60ir2b2xugE4ma7
Eg9MU4pnAUb9rqK+BYskqt2+YvBYBG4CkV3BUE2e27SAPRcTW29bOB8ftBB6hiVB
ipkL1sKxoZEzcfRV/Fa2nxv4xXCg3xPw99EVezN4AnnNGJY0WeFAeOnbLIaYT3HY
lBPBcWtPIUFrcQZAy9Hl5gBviROVWKfPmvL/XGFoZ286ZgwtSlh+GoKatu1ANx/+
2cgALIII1V1TBm9fOXsxb+8Dp+5bKz3tshKQn2tjgAiqp/anUXh+ziVmvLW9Nw4X
k3XnfUM7hiqkHYDUkr6k9JkkxZ32In2kVz7PCg89iaGEjdFVbenx2NPODtkOg8kE
RoSry8UXk1jvxoqXOsQqfKwmY6mG+k4tOH3YmdHsMNvzYwbzbN0KOhvozVBXZEv8
ENTvud35wNCe77ZOpQqDhfouIEbANZt10l/xqDHWUiV3ikZpOFkdhQPv4GU82VYk
cDH/YoHv+cFFspUniryGQ08ro6Jgp8wHfJ+YSJqYxGkXnayvBa3eeh/Zv+TmbSrM
7FDHu8OBi6NszIDLyo6vaDiCkIHHydpro8XvH0cysoYNTYpKQM8f2Fk/UE9GgAb+
45qH+rlffSYwLDGYxnAzirV3095B1lLL1MiwmJYYKM4O0iZHLKFe4Z3dqe1Ruro5
3HK9zikGHUziKnGCVGafmrZUoJsJ513vSoXmo25oiqdFydaILRpglVWMw2lqvvOk
rUqt7RWXZYHxY7IrFDhe4xzb5w3IMsDhWC2EulROgsarIcsmenRPcHqhKrpyvFT1
w9imS6VxFuo6OSp7txrdfgN/WUY4btLbf+Cc5cVwugLYVPLpf5U+IoPSCKiSCaBN
cHsOqHpvvqJL9GaFcEX+CusbSXSxrCeblilZFAT94RKtg61dvDV20HPSZMNE8GpJ
Dl4mKSKG1CsuPuGNZJRfXi9+AkYm687juloS7F0pSdazXSKi6wut/TDdNqTTWwTx
7svPELk3Z7tQdNJorSnKufbjP5fsNWh/RtokVrZoiCD+cduTWpzUwIfJLx10XYw4
27m5MmAIJe/BF9zeqd6tQfxp10ced9GmRsqQTku3AT0MBo/5clItDw+M5wOBSfCx
DJQJGvgpSVU/PGVkdI5JsrbgDG7z9Ehgz5W7nQonZ9Au1sssjTnQPq/PI2GPHBlT
45AH7GKdTOvy2fOJBquzjIZK77lPe3/Q5rajzxU+MXolPO+LTzymT2XPH3g38J3b
CUO0B29f54LpLIXdbLCoVRnMhm3UXEVBNwVCJ+xwJb3AkYvZvFjTKCuE1UGTHxv1
E0KPFKAdxoAgdeMgESNp9XWpJ0RD9MfbdwxFxiAbrVVQMr7c49fuB/w0q9oEKFfs
N43QSKEXDUf9Q67wyH3eEmMP2Q3YQO+kWXyRiiqlJZgGBMQlfgc8tQmNqYLAbRu/
U+HBFJe7YlFIinVR60oYEpQBMeTUt+2Oflkpi/YabmT/McMnzNzldB/2IyidVAk0
rso3fSDwDs+eox1kXUOqgRP0Wndt51Y8vfk3RyhTIZ5lzEa50sDzlpKMJQX8Ajfo
y1VtBFaq0DXEFJfnfB8punQp3ymB1h9fs+bsYIM6SIUgA1o+eU1iytiDoYL/L5+Q
nNwsEsnE0RijdmU8EZ1920mCLYPcO/umHzTNzR2nN0VOMLZu3SqUmkl4wtj/ABZu
jKBA+UKqePdJz3mndh7wHqqmP2h9s+JglgIf/QV1vD4lw2GDsnShqwJ5JyB07pFO
KQn+8E6wBubCst0ZDxOXo9jWer8+P0ME+qPZBdMuXo3GQaEDEgjXjrXG01ZwWLfv
YLSpDHrAz/KoryWxZqrvs4SksVC/Fx1FsYZQnVOLQooWgMSucYW7EGUaitGTQJ96
3bIjP6kTT4F/iC9z8riKPCbEE2jfq+MBXz0CcCBIkD6Vztqqig37H0mkhtbMZ05R
OYIaW+WQ7Hot6vEa4bhk2kO3bfTdX1EhpPtuncH+9WkD0ot+V8f5kNZBz/jlQRLR
aUTKtEZ9wJsKPurv8S1+wtq9HmXvwN/BpM+xKUrRQOjFRYk5Fh1msJUv8CA2y/PT
bBui+R5xeHSBgukthzfnybyUFqJ3YVZ24l99UH8HvCS3f/f/cIc3ODVllr2xeTyc
z8wzWtmd++S9Ctn6IXDgPl1n8SwKbUxfZYhbpOe5ChCcy9UR69DKZ5gEJ5sJv96P
gmu4OPmuFWDpFnkYgOCS4tVFlJiOG/3tx/6hjbuVQXVdetLDo2AmYUVj1OSU9wFV
Rn3cI6b7Xg4llKh8/mBPfp8ZRZfpQ5ak/WaZt+DnMW+QjgGS5kc0RqADnWaP9vZS
bsZEY8ddvGAe9wwt3ujp1oW3Jbs3OXPjHxBaYRhJowkahBELE7PS+5wiJcgnvNZE
b2WO9ybyKqUnVLemj4ltpP1i1r8naHtRVGNNJdJsQXi1OPW1iGpkPnjy66uQ9Vid
sqi83JQqIODsV7Qd9h2kt/RvNWtuxGDJENctU+mSz1LvZZdLc7CTNjMnUNIPgAtb
ymXAfgbUjC18poQqTpiz5iinKP72f3tIA25FZLZRkHkQ2TwSjSJzDAondWTro6ou
5GTsgsQazOKyqjvQOH4nMqrIbndRxVkIFzKQkvqR6E+1smj7MGWEDHee42WZWA/C
hBYlCU0KPUtbi9D8HPlvbUD9lb70lXY8+mdMdq6lzzCTgfHUcfnDhfwoGurMtHte
by4ZSkRPXNxXZWcKQBRTax7lsMoTXdmjTA2Wb1I2t2k6gMHcAS4/6KMa16DK+Rt9
m4j/poR3gpdr0BiDEjC+I3ZdYpEijo+eHAHy/g9RRYmKM8l0s8lJPhT6V7yfNbo6
uE2lUO2GYSw0oCA18NSmtAZk7bITsiIYSftWWrITmQZqVNJQGKn4cgGI2G7IOEI6
wZMxZVoyFXIYUQUWx9xvBLVco6R8zGDEjbwpgHWHGYtI/jPv/nePJssPbrvk6Jij
uffWc+bIJvGHQNI7NpCQO7NlMwKt9oLSGLo+Q5ML0NIm9AH5NCVRAQlHQl1m3Zn/
w8AyqwPfTmF2AHwi8E2gfhd/ciQwyCxbqFTvmqCZJ7mQQuNSOf2aB650MTNqPkVJ
QGisEwEmeKlocPelNXd+OI/2V60MdXh+h0AM7alm79bQR4VuekAKBzCbvDG5RlSX
2BfoThRp5O8E3qqGTljseN60VG193zL1l8NCkSMERdFP0pEL0L1KebdqDfxdi3lE
JDqVSflph1fCG0zBnrmEBLwEcc9Xn7aQH+7z0jb8uao6WIag+PWDUAIhPnuCzxlF
doEi4lM3cqiwR6TGZC2TRp32NnI75TnUdHOjCCsY2LRQUgfVwou1wF/Nl1sXBrsS
9x7qiM7XRkTBirLEGgA6us5hMbUuVGjA0QycQNx8qSuKDb/CDHhxnJJjCjTfjmlR
X4xHpTniDJ0xZZnWKBDc6ZeQ2IOjBdXdmkMySwq/CM2kXPXADXzOZL6pPcwVYp2Y
O0NhzfyrG4rb5xuKtxuIcjcIr7niCeUSLfDLU9EcW29wvOcxSnWwLdmJqp/U/pRI
MJlerNq6qm8NoqN0B8TDqPva54johsyrh0rBrZPEFAvoE7UC+w26W51Ya8uB1+xW
CabHYrReqLwIScyl+jeuJXVoChDgXrL18sdLATJbFPOvC7oW+mRLapU05kEDhOhc
mNPW86DZXerx2oUrKgf4dhunE8zfwvjc4nthdNB0ZyUWiweDDeeY6xIclxe34QOv
ZqVz8wsXBrStYguMYEAbZT39nCVlOVLWdctv8719GDPFKtWXhkhkvr5HgvONaxuK
NwMifrD7KiHqQkdi2PhegOjWbBjCd2Xa5f1paZ/+Gw7MJ1lPbXWqI7yi1I1giSBm
8c/qkUaPnw+I1kUxa/FDWOTtWGAsfU5GJEb6nVaQv8CNd3ewaHflUY65GjdQ2J0Q
09dcO//N41U0DdvQKlJ4ypGEc6d85LrK5UCtD2TK0aVGe9GsQz6NzXs1ZvO0Ge0H
ekH43m5hsHvjNEL3S9zKFJbRBHlgvgHZEAXqIeAOfmp0HzkPCxzdbiXMtTNOOg5i
Us5QgrXcEjcgq0ursLBWn4GOOH/35QRGC6/nwj70fj2i1QT92UdrOBPajU5ulhMk
/F1arYOx2Dv2rbqaHFZi0feTUBuO42IFrtjHS03ACL4Mxw5eFKrgkcwLZVKguzuZ
+AL4ojeqZ6cbqx2Ra/8Feau7MsGPFgDbYsKM9q41bvMsZ1bhXRaUZyKovGhaDKMD
6+gkFHqABb26mZNN9EXI6sRzShDIsKOxxuTGANPGphJc9NirLQp6UTZKzbmc2e6z
tywDK3TtoYdOqFFZvEjDjWn2rS3WKCBoUfxsn0p5lD3CwXjONmxRaCbTFHxqomAt
g9tyrze+nLs3lH5YH/pI6MJajRBsRe9gPEyDVSSWDKTK7TyIrhPaNnwtk+qDP2bE
6tusUvYtIMdmsCs3pRQVJqfppVioG2KgKnjYpcQfd5VYGimChcuReoIAM5JD7CnO
lW0gdtA5BwnM3p13j/UwHpSwd9/dcHb1a4RFjaXqX6IqEHvfcmykUCNA/fm+fCT1
lywloSHiUNvuD45/rk8lm+oRw9UwPkia7Xx8I1197CqPKPRydUPlSVntSnp79KWK
WXPMTXNZrj9TtHGhI5OP65IBQkM2x/ZdjiShPhsB7VypUFwKNdHS2pCvcFGFpn/u
kR/YiAv1MkfxdGJ9yJdOQyArTDi4Tc8JyJ3JinJB4bME6vMcvshzTf5g3WJserKY
/9FVfkLS+xQk4I/ydifwSGlXNMKLuntPDe+k9+EARG+SUwT2pEASrJE1mh1SOJX4
0A0JklD95UGYM6qFpsA/8bzNdbuwWLim1DNj9U1z7oCRYcxgyVL55aIXkAXzm02b
zONP2cilHbRPhNhWIji4qp5mKCesFieg8dgpBnz7/5ar8F5AbE9omMFk7cBbPEYD
8/qtTVnT10cQP2wT/K5cwSWvrL0Oqpxso0SYmDC04r+prP7mOoymgqmLDAWJNXIP
EAi2VaXFyBKtO7t90VkukF/NVbDnk67Ybve9HVaXJ/V0ONbGLIXvsV3yUasO1VCO
bx/jzQ6XkXyPWd7QlhuLVE0PM1TCYJdNOJNJsQ1gBYEcAzMFdE9aqOq7GNtwybfi
qxqe2R0NfjR52Ecp+jhpXtY6Jl5/VPILuB89vONbvPG31Qvf0Z+80HhhOEoiBROi
MzmXr7XzH71Wwb54pAF3xWSLTzAU8prKFBKpZcFKfEBW0LcoYKq89qZSpaXJXnO7
FYk4PBYYryAdquOlqd+cRG9RW+uSywBqTbDEoCMiVxSHQ8qUZTxv7BrzYct+jdoe
/2qo6Z6CP8eOLiEb9fVdzw8cIQGsIcQTGzKhEELHhdyVCmdbWqZ8y1VclHkaVDjo
4yrvo8XlWnRq+I6IOnW/fnkupHIJP8OAT02u8oddc+14eEapRlLJU9Wj0ee66KZ9
EHPKulORF7pCm28scg0rfO0SjfHUl2M077KfzaBf2RUVuUJ4Z2YpPfGQ2dGWVYLM
o8FqWIl1AwsPpDk+ovSo3+iVcRo8KWmd4ZzEtcQF8G1TE6PeUxhbv0KhZYKtxtZD
wLW4cK3swwNAoN9IvqvCPvKLz0bhQdvn1DESRoZVokozfDXsunolk6FRmplaE/MT
w3ZM2HUF/GRhYUbleHVqeqFMsym0DcejYdDHxhF0zIH2F2SfzqIe+TNTEPWQkVLf
n6xrMWI7yyw6eSWx7p19tzk8UGTruUZNDxgmunaoYXRXT22hBcgq/jtwnmPMzyuA
YIt+RN8BvwoUdXJ99GheHwH4fkAOQQBFmlOxeU6DuoNJK6coVIEDfwQLieyoQdVT
XREg5yvdjQizpm2FrZU7ZuXbBrWtpfO2bIWelnRPzUBeyRyuZbdOV5N03LL38TZi
Wv8CNZVTD1Dz7wQEy6kqOi4fauiO9xe9CHSgidXw3r9LwyDVmFF/RsXBUnRgQcAQ
DNokkSyQaJRYZV7QTvAr7lMppYNNEEHLxu+A3HRPgCuAvBnHJQdsHi2JbodUsva/
A7rYaphCr3OmUOSC7ccyUMXp2PMzp6u6IE0uqZqlkIVYWsFaEWnEl9GW90ACignI
b6ymBSzfjE67C9fDxyWSSs/rem0WMUwGFk+NxHjZO42m9vldTSXO+OP5kCDwiYKt
9f25MZi3XczlrrNFX/b5vqAz8XeQ/6gE7qnDUf/K3ZBTDuf/9D3M2+B/frnxJqfb
BvksIdZJrif+cp3z3NKVCkwXimucHPgFY+HVnm4eRTwI9jALUIudsfYij0cqhvQJ
pB14K9HOb5BcP1UX7qm77m04vTE0Jl3rOPEoeOF0Us0VDUhzGwvk85bLh69bNoHI
UuMi8zBN4bGI3mTB8PTT7+raBY8qrGETgnZlky6HTHNXzrA24ah7PDkHXaI6e6n1
cYwP8+31gmF3srmKkjI2S7/Ofc43a+di9puBqhQAI0w8jGVtXRlfGachNF/cdcro
MpyXk1rSnE+ZtdsATfNr4O3s6VuC2554+b3kUn4lq27vPTVOWs1OrT2yF0hkhSh3
j4qwQmOCb5Sh74Imi/S9Iib06IhGJwri5FW3bdoDl52VleEHOrDy9cEna7PYiAnQ
W/s/I4TqyafaRFQ7Qmd5obb30NFqmcl9+cVZpYFPQoddtcQ+Ez/R7xyjQZL7AnN0
Ri0t2noQ/rBKk0yJ5uWUqebrFq/EnFyKNbQPYinJtZ0UKtm82p/mStAiqOrHNp1d
pCpeAYOQ2g5XE+YYILoimwWii6yBIQyjFW2BZSt+Fcei84+R1go8MlHI3M29Ssfk
+jLGDk2YWw051RMDaJNTBwv6HrfIOEcWL686NOy4JuOGc7Y3dp7RL1QUz6RyQOcR
9IlRTLGt1p7FY3olFTmWZxozCRExuid5iZ9OlMy9LQb2jiGISwzu0oMEWg5T7qXv
681+rjchooigvi5k54jkVPqYp4bfX9CJqJzJ5LMq1wUX5ExKwKy3EjXwav3GjcXf
rZGSLJbmWaE4uXxD2gpGHxKVNmGfkJBdVBJekPPR9V7D7TCLzjnBjZLCAakxIp0u
tmXE5cqIAk/u2lMv/chAa57achauGK5paPxnsUOr+WlZPJ2XxTgDc20kMeAxRDM9
EexHHefGN3Dvtb8p9ZTclkDdnahCPH7VXttPujjD1JrvUX1jCC3EP/hWHhVuTbrm
rUaey+BDbO3lvSH6q7ZUFg4gpcK7XuDzPhXng8yKgBF7e5IIKFy5K5L8ktfYSsbJ
JLNqy2GFYteFQerfYMV1p6vMMaWCifaQTVcIbGXr3Wymw15q0wVCY4+q2E//O5gg
iV/790/47LOmpZBHEmN0yb5n/peE+rRx6Il7ixZrmYe2QXT9O5O7wNj35aTcefes
vNwtR/rPYY2Oz1YRozMQ3vyobv57Mspr9yNa8l/DXgx779cAJwQZbIEV3zlXI7/D
tD+hkrCBKz5f9FyVd7Qox/IS782WKVyWHkV1MZCzzs0NkJE+/0qhVVb5QJN12YVB
EGLpc5k+PDZDJcQscIOHWODApHmyBSNXnrsYiSknWGbC7QZcLCwsJovBU4/uD5R/
bIEMxzly5rtJEMoeO4ZyeVK+EFMHVQJDgmLdPUZ2lyWbLpj7uWwY/rj1XMvsTLn5
KTkc++QS7w5KqHvJ9PjG0++wGOu2ivfSZzYpKiGOd+26k0/d1gS+PDUQ4WedFtEp
X01Eyo8yDZpKZ0JkCftb1b339JSDmlgaaE59GsGv9fdwfJQmp4qznatqH/trhWwX
bLEg7f2Lm9wcgD/i4G4wqvlh406+/CYlp3507/fyZahX53p6OUxExO+g1XFZqP91
3S0Mddv5FxYqBU30AO8UY/3lzOLc3MVRvNfDo9WjQ+WS14WlNwIN33rH3nXx6Vhf
qYDj5ZIIn/rq6VbweB1moZCkoVYsFOb1D+mh84OEYz94H4PWeRLNDj+uHec/7+GQ
HyVKbZ1ZDk7LnjK/dybzoKO7EE2LYDUbijA1nqQXQjaiMCO/F02A9K+Zitmebt1N
K96F0CUIhdjMcUDTa9qGk3j8oubJaO0DzG7gRTFzqsJ7HjpsZt32qGa0rAkTYXVU
jflM6pAbsBewhptdRUziFHAg6WRIOTpIBMH1XpvLPe9kh+UdkchXcaMHtvomfRUA
/LftLSNubXjO9Jp0P6YDlANX8hYUlI2ZqB2xhFT5ZirRx7t2uM1x2ZGG23U5SmR3
1ax1i/UcsfH8WrDbA5xfC0Hp2fd4jgc1ne585d22Z4s+bXnMWFG3sgRI8IraN9R7
fIGIDMR5X5hj2Tw14pAIx44tawD18oi7GBsfR9e/5+pgA+tgu914DNRoDRx5iACK
6tnuLYBfbDf+Wbf6IJhRs3JHwOApVGOsWjYpfuJdwMkjHynPbNokBDoUS8vIFBwt
3FijtjTS5tuGhz41MAIaqrepU7Hmdz9qFUX+lyR+2bKgmL67DS+y/lldyn3gEFVZ
si7x1L7vj1+ey2vh5Xs8ZpVKHgDI5jxNUO2Nmr+YmVEFv4BLWUL7NOh3Ygh51xn9
GFv5/Ilre5wgmUT2W/p89wNfhJCBKBWptd26vGxFnHuIXovbaBMr6h3PmE6Nv2pn
6T8HaK3OM+LN9q2pcS5LQGbEi7kvJNV+F7TOhIzDgec4AKEatiGibBSCgInFiZJH
ikC7AQP8h5lNukgH9HQKV9L2kDvNA2OnvVCG1vLWUjLoLqLyYE9GhJFWhw9Gewn7
HgCu7pl4700qvN24iRAYA77r+Ummmba/FsdLtOrVHDMLyp9yQl1VxDlRVL9MXAM2
ODBmfKX0z75dbeccdy9XL5jDl93EmCbYkeiHq7uD46qGuF6gdRPZDg0JftAD13IS
OlX0XJl4kIQuCHwgNI6221TJdxgm5yv9pC44Fi0oPwUFP5Gb4RJi0J8iAojM2/TR
RnRWuXX8X0D0mLCOKEoOxLqmIJfaWInUT3vE9gLcMGdMCnW5IxjvMx+FE7Y+xwRe
iVvJ58ZfBGRWHWtHGgrH19KBMwnlYmx2VgAHnS6Uira19/j65PAUHCPTg1mZwY1N
WQj5ioRn46zn2FzsbvF4sFrdJDWIEOsV5tNKDIDCgFmqabpa49R01iCgsD9VRg/B
8rMobYc1NoElnI/LyldfaL6JfpqDCPMw5JruCI6HzqKPsF1sfniKl3Pmu+3HY31/
UFxjcA/v9O4GJ5hepgdmPk7LR6zN9I1qizBKyBq7ZBDscXz1uSinc68oy81sd+pQ
gI5KiavYOszxQq0nM09oByLsmmGWWSRYrmM4HnEvdZvhVx847676FzwogAjNyO0Z
3oXgtG9VDrkNS4SI6NBFzXq5D5dkgyGHKgLHzL7+uqmcFRhZeH9CKbnkqZgIDInE
lKTUSRngWPJZDbBmLCeq4uJIQHhhv2+cRliNHl6GAkwJa3QTY8OES42Uij849NHB
O3O5FLmJtMnAyRYvW/nVAc65uijw8geVQdZiQJqAr8LBArq8TOuEcbODnBdc1cSf
gTkBYepLjvmRfI7qDo3XS2fW+6tqTdZ7fHEK3ARuar49iF0dp5vpN5mcfFD1231n
L8wWbtrPwjk2wc2MIefj3wjMdTL66bhHXIteE9Cv5qoHoa+YQvZRnrSYrNrsTzyn
F/wOpX/sooNVY9foF5BSBa7GN2sfATlztuwP1hnp5k1H4NtfezbHRTB40ZqoEt5t
1zZnerJfK42uLohMJyOYCuYQC+BWXXPAUJs7MaOK+3nHcfKRkCVy3U7b4f83kAW+
YOksjJ63WkZPS01MwM9AL5ADJejdilGh4E2sOQXl1TxeK/ngFCuoxSHn2q7hypug
4kyih6sc0MPVRgzQqkKICVJjCuh3k/YZNUuQTl/CiIE11uoyheNyFdWiobmRRq3I
IIRR3aok5xO4859OFGvIyJhD1Bn/uz7EhENjwNQm+7jSjx3aDmPS4gqK0Ik12kU8
Vg0Zn6mEoylqpLG8bHb6mpkJt7M3cUyYtvgJni33hdkEFrOrFzZS1T3+oeX59HZh
Hfb+eYKQg9ATyCg0erZkmivImOUaricB2NCHNYOG1ux5tm9d8pI8bjueYbpTtEye
ynV7IRYxZNZFbeiB97JYYu0ilH6muqSGZ6DTJVkgb/w+CeEjESae6dODNl2/Wr3J
nNUdjzmkbJR8YC+xPSFziqofdMweE/xkOr8AS8blCe7Af0Pon+ckoEofCV0xAvqG
QXdS3O9dzdseXbHFsHPrUxQO4iUkjXPGf/EEFBjQWfO9HvbJMCQJgUgZHvb8AeQC
yCLmmOaj7mwFpTS6FpX1ONEJ2r57bUjhFP7vAzjC9v9VNybsRi+6ZSCXXObZ+cWg
UaVryCnOa8lmR6QNnLmal8QINV/7tVZsTsERV8Wt4uJ1di1nIF+XZzXr3nB+2Oc9
Dott5rjJrAQWQixoLCsa1lThFlcKVlUoE3/4ww3KEnHDzs8oDC0HCVDNI//AC71d
gNXyyg2/cVDXoPw6tlEBI57Au1IOkiBslKf7gPbM5/HLpYoi9HDsu5BCE/Ncc3H3
gAhH2VqJrDPspRIffqa32thp8vzddZa0rRSmHjhsjnrs1PzUltS32cigZCXhslkN
KKn4PyGX62FZsa40hVjaGYPuJEXSz4AWStJhQ3dBYBrhUYhZ6yuSEsVvkXbRTYoN
rhKf8zBCpewOkVz1N+HbqYs4HEv01rvbP9S9w2a209+0aQFF+VHcpEgBGjfmpYDB
yUi6SQytwjQbvO9RjZUOqY8VvwY4WLFNLDPygxiCjqd0JiFjcJwUZrWzq7j/xaLl
9t7swsFfHxuHHzfiFeHJmx2proJwpESqlSdI1V2erdt7kZMkGyRq4EGPuWMcgM6L
UjJ2PsUvMxyWAgzq9okrHFudjI0xiMa20lWcnYB1FKEySbxJfM5YA/SGvYvMnyy0
s8WbFmqfx4nqaqvf7fL3tICG6Rt1VLxJanCPImU59CCbPXzH8KJeu93x6RWTjcTV
Ee9izJvVIGB8dFKYVgcLPPSyDcUgkKu45XH1n5e2zdIiR8BMmgqRGLgFD0hwiJT2
ylSf7Ixpxe3fs5PHxrebU4vobwnFOk7JzPat5cupiGUJZpZTEY6OAsGBoXyAhn8Q
5hm1j+ssjoD+TEqYGcH729GeZ+03x6qpWc3Vd0/QdPrXOKkRyjhujtv4ugxDENcb
xnAUdlh58Ss7h9PbdEs70haIBi13GUzr+uNgkhnFHfBsh2sEdPH1agRaTionLEsg
kV97rkPZ4PBbA+jAf6sbv0rCWjCoZ5foemJurZ3LG/tLfPmfb0xzIQt9+UaIea/l
wWzxfCmxuJYzRMdPTA5iSP/cr7LaKnjddcrjF+ZCpr3CoQo8L1PwhTaDvELhbCef
KeNDDGc95iwUAPl+Sa7eXjRSuMaOveJv3fx0hzxpatMTxU42TH0C7eSiMbdb6hkO
ZWtSgFF+mDjZnBf9fxvR0N+ScHYp0Hz8UgDhlHWlozJ7/ttW0472q/RcABRPAZZK
UlkQDJeBO88wOemMgHRx4fv7c1rRfX42Kuv3ZSxvw9JHrq0mLITpKwLYyPLdPDia
j0tOEdOm416+TCMeJVLbOjxMnj/kXTYxB3/0s0NhExSLnRaXo5CxXPDs/QLRgD+u
Ais/g4u4e+KpNoz7dM7Lrlx73uOx4PwpAdArghUwy+1QHXGuTP5pfqaviAi7Xo7G
viHscLkveGqDrB+Epbtr/4m7p9iwBfjHldxuX7sS/Fp15z0xlXkqWy5vdrxTX7lF
X/ma24th4W1g2intcqPN2xmoq8N4+gEeStSGWvjInn5SQt1eJwcCMawXn2/QiK//
0+jMXbo2S5lNzNyKuf1xk1bYX+YE65dWkn3Z9YTYerlj2+8XGrT4RdY7Z2oZOnHn
til/GIu/Y97zt7RoH8cWyICW9kxXkbpjn2dD8uy6Ap2IQvhIUURDqnQM2GhDnBkW
OVa0PE0qeOeIy+ktmpLse24uMuAvyWkpZweM+7yvj/KI4AusspXzMddxkakrb2ov
t7zZLiHyrxGTnLRwD+WHE4akD2TQO3u0ltAzAZ66LDFaZFJSr5RWG+s6JjkiAWxa
XHjZV2n64aDBq9pGKgNm33THZ8Zf524iZfWo/9dVENSMOsWlB6NswHm7UopJ9Kzo
+4j0VWqkB+S0jr88CCX+tXd9Qw47XiZltLHKe7DfkbY0tzSX9k0ofOs6q+5HwHZf
GsviyXjALjsYP2vbhxZ0Kiq0dNPkdJ/haruGr3HLuru4afcZOQCYvX+QHCbrSXsv
Io5p/SyA6klQF8bBLoX3W5hOmmK42od5RX8y8eXeZ2SR8cKI4725Oq4t98d8Utb3
L4ZfNVDuHO7IbXG0sPNsphplQAXz2oD5tbZ51SdaJWOlWQd3+fgyAvhpkzrLW53R
3wYthTjT5jofi6YMtrhxmvtUModEkaha8hSjB8+TbdFQJDeRY2/EKGuxrxcjRWF8
oa2E12V8+j85Sk+DPlq6OJmgDp/Hz92hNaaKupdjNezmvwPg35cAMffSlHps1a3v
5gwYypCWmVbVBLCHbKsXz9FaY4lx80djzYbG8eQ/oC9rRzwp+QcjtvJj2UxFwvUg
iIC73DDZXGE/FR+DqaAWKCWwlAj8JbSzF1iJe8c7w6eZGRG9Xhypth50j80zcpJF
OGuTMJZJwpdAnZizrVRwd5v/WWWkYG43MLCDmSBXvP6gQ2Sm7T378Awp2JMKoDYd
AUWIKxNR9Tg97nISYnE/j967c7mpcKttfIiOKJdvhA8aOcinqmfl9HH0ef/TRM+J
bAVk14+hPmGIfrX7/J7muncI3lsef2/fZWpVvqSOfoGPThWrqI5D0USuV8cDbZ1n
iYXPM/VoFxUdsSDrM1rcHJVb7K/CPNrwXvFrb6wjarjhLywelGQPbVeHLTBFSIyg
5AgW1o8a6DjMO2BhogB2v2tSNts2saOAY/3HRrHS7uL6pmPwF3deXf2pa0lFplKN
NaG0CaXxUP8wBYbrbmENMCtyKxO4V8wB7OEbot3vJmdANHiGQIjdlQVBoL5sCaGp
VoiRh4yZwMj/B9ghIUmKWj1E6UlWXhGpS42uQxZxB6vBgOiceWTG/KZF8BZ5g8Pf
n6fFGargDELvAhRGYmUHOvCrq7r9p5PnjUC29a01Kh2zkAN36BoDvvC0+mvD0SIP
JYJnj0aqWmi73zYftyVNavkWcrRk6xPzdB4Alv8Jz4XOHrmu72Jv79jqEdQXckL4
wXcTfj4Xw/4B1msHiU6g+kgT5tMl3aQgsWseLDUqDRD+bD/EXQ+43C22nKe15qxN
ZeyaN8C8CtDaDuDT7kolsaL1RTgo7+n2YkAQAM0v9PW3VFSZ+el150cvY6dOiIYq
AuXLaBBQ+2X7cmP92k3w09x7f/iQkULek0X+DT9dpA96Ow99lZ7wGl3Jrv1y8Kin
gANiBeHeqwbYDYE6ZszMnc7oPCCjZW168qfCqpmSREvyhv9JXXtv7FQfWKuc2q2P
fJRfPsY225QY1OghTD661u73gJu/ycNEdADtFe9TUSWxmoG3t1q/H4nB2n38eBly
vsiM1yqpXQQFF26UilTB07w8B9Yqnbxm0J8ijv82ueWV5/k3ExWGBgLixzFBGUwW
AYcwOxF0D/mfi+NQsiEKz30arEF8tMaxaRYRtBw8sRuG1+NTO8k0TI0NhFfK6Qrt
oFug1k+5DqMlS9ctWsM4EjZs3RHTWZGnXMLMNDXU1Smb+AWz8aqYYC20Y6nmdeId
KL7Pj/nBQFnWZITh7d/11/OU+IoAgmX+klc+frQEMX6OW0h1MA/UpkV5IFsjwbNI
vuH3F0yuFaEyLdtc6S7hjxkqG7H4Smr0nX9cOxcbN7pQgWalnfS9m51H7qVA1qcm
3lxakgdBZm+iAEnQiZG3ScynzrWIKDDk72eGQWQ+0nYvK9baRnlDXNvYmQaB1Qu9
HgHdhSkcor502Lxaq7J7z5cHMBekuKsCin+tA3+ytIx0O0EdnQ9YlFDFVfPJio28
mmvHWlEYLk2Nlz/MxWXYV10Sk0fgeWO0YddWUy+/ZOxbG5HwpybeVjNPBdIm8kU+
q/uyNKEZlWJh1bjEW5qqKtdo01y2Efj0cmVzQdskjyZmkrw0bsq/4eDgi8fN/qea
XeyUopWhd9f6sv/V+4Ch/RC6BtSYnXEyIUKqx0MQu8EKKz0hMsrZXnpljd7kLrX9
9zEl5Zz3cAC2m5TfGUpaKukR8Etpx6lVtc/isizx1QkasoTgtPgAWwK7OSKCMZQF
jv/uI6pLCZmktCZTZ0gbNP9mcBJdmqyJFKj/RGnmmuTrBa7nz2YBAJQOX41PX0Zi
x5ULrDR7NXz9600ciObCdy+xSqV0NeRhEqwxLa9Pev+G8uREJaWs/Gjt5rBsdh2/
sVzuQ2L7IM1i+AuBvVdx/UNNXvbLE5gtm1XyRwxijilce31aMXF/dnhsY/yzdUCl
H1RCg1V2sMphwtBL4I4nZucP40kykBZAdlfHnadpBOvjIvMRUEiDe3UoLlrpyieI
eygeHzaz2rD6mjFKn8G253NtuZu0esWaZAKOvmes9idycY5UQSV+nuED9L1SVhMb
9Qnp8ihR9FS8kl20geI1Bg7EFRbUPVi/KpHzrWGS15agpQYy5ehMNPN93s8Z9FCv
XMPYLihixJLp1YbGzKLnWUu+CcgL9v9PT+u6UFsBP8I+XlWo8EjRaBmV0Yge3dyU
i49Qaimb2wNR8bo7MIeBpLJg6jLSatglrTXyJTJgb52lULVDoE9+tnIGZWsxVcMU
4JzQKt3oIum5NFtXNLyKYiL2gdjuY20zKsvwe2SIchs7yVQq1G2HNEFpuR5Wvv4s
6vQ59I6CFfkONUOTj6yC8XCIdjDG7N4dRAPubmlOYErYrZUs1BBr9stsih/DpBeC
OpC4Y5OPgYIVIEWiFxJYVmlc/oMU6I+QmS4a7OVTly5jTfUksFAwzvuKa5NpMCHK
0FPQWpPeJgyAO1b6VVhlzq/CjFrVTitQD752nDcOYuh5mhNjHKyrvibUvK9ae53E
cRhBjqJleco5VyOvumoN6bR92D1qLVGTNzNjYb7L8WCjdzUu9U5ZFLfCI7Oq8UOq
tUWCR+nMmW3UQsEWT7Lx8iUsdG9YvSGepsYHTt0vahHN7AOmWK81AXbmsev3o8Pf
rQVb/VGHljtJmMP55PUg6fVxnXUgJUShH2Y3htm+RxpopLPaOFpJV/zfOt03HKPZ
fm8GHXDbMBUZiyCjajuopVQ/GZWOWaVutrcEl6y9Z8o6/gE14OUZM1aqACjFhecW
SDV4bfjO8TC5E09NV0jz+uFWcFntSWQ1MS7AMaFjlsgSyiP6zFz1OMcGIK4zmLme
G/8TG5IAj2rVcnPjhzbcTF5UFoJUiWxHEMMpdbGL4M+8f/vyILV9S+fcomoOvPzS
wAHvbD2CU4PNSpTaTjeniugk0iNMkzKJ8gToptQHcdtt3bgkeIloJCdhjUfAti79
/cTxQmm7hguqLbyAD9wdGqIcai6hPQRgIEhOLlbSVNJi0wSX0mCux3mUMawa1z9x
EtDvcZUdafqZGcoj2lwl5uBlg5UPDwoGnmQQiBXQ0HbK/5vjFnEej/1Ee/4AirI3
KiRmi42uhPJF4RCoxTrrVDKT3TNHnCZedW5zAqphFHGTZMJLKk9MeQygFFGgtd9I
u7W8LM4naFhwrKT1DBQTYzI50xk6Vpa6UovAwUpLjuEptcUWJuVWdcQZ+8gqaCgM
SLkeA77p9gj4S9JcLTB4QckpGSLSKV+L/mfbAiPMK9yuYu65KTVDixGUeTZtOR/A
/66+I883ez9UM2FWO0uohXL7ozF2dBqqWbyz1xB9ezVPn9e1GnO/H9DKrMW6W7cX
wS5Dvi09XfrCVBnoeo7tbcsK5NpmClJplnNB5S2bVYID8T6fOvVKgkzSMFozlCxj
92jL/Mg8snmDGJ8Jsa06WIfrT3e+L8PDBXz15k2jA1TRiIxl68PQzs9gI8hZ9mAG
vajSEPcYhRAPc8bs+0oGk+YrQpNxZLBTQcL8/wbU+uXYMs/elVt3Zidz94EvBx89
Gny90Y8y3sDYMeFngEXrpmjR8Mb/hvJw4t9GldZdMp1nJc/IzmJ88PiT+nIDGFiQ
9HKt1PU4GFmQrzC8ZJjPj3KtBYXwqqQOzz2hdLOmJHidVe48QY4XRKEbqv2szzgd
hhUwOxGPLVoy/nEZrA6HajfUZcqUj06RGfs6z/hQcOn/72soqWl89NjKrGPdUrLM
NjZHl1MKdMV2SpF7nEbaSdPCY3thp6/AM+OKsEqkPMuqETWh1ETRzJjwELLZaFpK
1fJnU9/gBmL8cWahinT73fKQdNJC33m8Tly+9Tb03sn3lHDXcL3Kk9XK2hc0JmGw
UQx0l5b1uQ8H/QzcRlJ4j6vcr8DxqZGoz4wkZrReqRXpJyaURDbvwKK06svyzehE
r5G1lGvOeeMrXl5YeRv87npTc1Rmt+W09PDqVPC/Nta0mDvvPPpnY1De/fCX/za0
dpITNJepRk8WjkqDyByFsQVcm4cKNh7oJWmafK4Zk2WdNgsevqwV34sxxbxmSIUw
fgOIU+kvh5ER4pxWJLjXOiWMHNE6t5oznHrgsiPtO/XsIGXixxxMPxHyIdG6U56a
XBka+XCS90jsY3bvaxT5OtLkEt7Fg19y93Bsu8fVL58hJ0AgMiKaKjPCs0/k1HDP
7SDpF+Fizg/aj+00HB/KLzGopO75s2R1UFDvjKJQMMGgIR4r41XGpw9/OmXr3E/b
SGPsnmo40/yb32vADGrPiKW0RLwe0dAJymry3Ft48nBXqVZnCWdQ0p4QI3xzKna1
PVP0t4dXjKVq3SFYB1MDMaIjHYYXK1SzqqifMSulO/8NFkK+rh3vdA/+wzoHdpS0
uJC7beimutSce588DI7Cn0am3clIPet7UD/v24mSydmQ5J1FcSyGKUPtaFQAtmjR
n/I1Cy53r+WL11ys+BDFyO6pGwkF89iV3B9NVNp3oCLiEJqBHS0jdv76zo/MznPY
ejtxVFT75huGd+tJW4S0tCaWUMCC1dE+Gf+ZDf7fDdPSe8Mu/PDh9DX9q1FnV6tF
4Zs6MGrSdFelRZmc8QeOrkQpXkzweebbSLD1VOvQ+5N+eZYTXXOVq/WfQET87TG+
9UstoFu/AInTbiOyUDlGkhjx4/e5vJZYyYWMXytNbtQReoBmd1nFWWj3MmaOwRCn
XcferONWsY3xyigJoJhCVqfafm1NUKq+KXoETr0x0YY/tLRuCv68rhCyoPBP5SMk
MnacuDKoJTAFDU/8oIcMzm39ux9EOvPoIc1WVcBmlIYDZn4InUHE1NBZ4jLQh09o
QiheFwQeUQO5QgeUpp/YZGYaGSyuta7cpTF/H6oxsZJn9sl94/nZxprfyQWze1vZ
fiYymB26U3TJc+ZzcuyhN8kFXIpozsr2uB1My9hhL2iWgzrrDyKce8iIZZuVYDiT
7TaP81PE4QL6I80zwG1Dky98mY26m8PSycBN60p4h31V0YJ0VHvEUGbPbvC7GzAM
4IxjKTfJGJvj7eCweYboDwU0rEbujNVqPhhXEEYKYf77XRcloMuTWrfCPCS/8AkF
I1WWwA8QpDqcaK7fRXT/ezCtxXewB0qCiarNp92aPWAcTYzrpYSVdx4RcBLeYxxI
3sC5EmBaLfi00XwIPZXkBnNSjYXevbk/7ePYcQ9lTewaNYnzgH3KwpM/yymG9q+J
R+MDTJVPaQ8kk3F4Vh7WHd8SZmVUI9RaRjn366LmjrvPSBGJjVh4iecBTY+7gx5D
SKH/EHKaJ+mJBA6jjh+5p7oM22n+r3OhwCWyiYtY05/B0GRE8bHD8E6o7XHeJuGF
d05hu8teEj86k9htMUdKAG4rC2zcBvjxrIaIwxNS9Jyh/TPGcmRsHl8//M46PtAf
zRiyZxc1+t6R9FlKcLnqmtK4ZlohCtF8yijOl2p4wOTUqPXbvlFPhNjMBz4igsVo
FzZWrpD6mXHE3oHwP4wDprnQwVWJqV7k55OsIAVYF4/NPn7Xmi1FNbwCenR5nwVZ
QMWUpQ7byRbp3a9aUYj+qr2ZTC3Kw33UsH//0sjLA7FIB1f47NG00H4mP94s0gYq
p+uduf5mV0GSd2CWmVpGi6qbZgk/2QoM0qxGtwix6//5DQqzVbmJd/jJUKTJUEfx
lddhfW9PEghJzmtOdPDreYmVGlhtFOThNdeMTnyhIGwbCEih2/9rDeHd9fOS0/T+
9OiyY7wZpeD4Tb5D7aUw9Okvf5Kpq6zuo5lEBw99KnGgkfI6ReMvSMbkKBsybArX
Qs8ypBRhcSde3uVpikPsC6IJ37tZh3VHNqkKfSyHk29UOJd3QYagByEDwfmUvimY
Jj22ZtUAthrDCxqWrRVnuQtziN3PPrTw2zGp7QREB1yI6wuhMnPwb4KIBWgcMZkk
q03QXTfaJCB+Lk3PM6BgYV5ACmT7UqvKNAOWQdVRm1LG9NZDc/7s8i1GePJMJO69
VFOT0s1YsY8qlqADwvCA93aEw+6U65GwL3teEkQk8rNR5fWImsV8f7zHxRQ4DNDP
6Gc4RzGQvnAgUKFaQ+V+53NJ+P0y4Nf9ux2A9kYJf++32HAkz72yrqBDHTovJDXh
mD88tiAn3wtKSnuLuOHIOCS6ssxiM/L39OYBcLiYzlXjtsDt1cw7691fzJ60uX/x
kI8/5n3x6x3hGTdmbQuxRGNOxqARpOc6Yjm2n93QBBr8fAq8G/S3g6l6i1yP0L0T
0gT746F7O9qG+g/gC5AZXS0wPtKOjOmnRO8sJF8na4tQillS+89frs2CaaQX0L5C
4Vb88Qd9+efO9x6lhJ4/F6TeyCJj2fHNMJazuKi56hiDchTV6o3nkaZACtOn04Ds
va3I/kaadePK3+IUVRusJ4uUFCNGPQ/sjVcchGxzq088kXi4nSx/EU3q0EH7jXBB
QnhIyCFJqgsFq82rzikOFdIBXPOFOfHwC5NELD3S6Mw3KhvE7b7Nm38tZP7AOXlr
UxPOigZ0ViFG4Ck7xPg4M0Anzypl9KkZEEYB49pAfyBSwHkHmTgGSN0DsWSkO6vS
ydnVMlEH1KnKH7jnEAuvhM1pr4xtpvCvXqTbY+LOP1o+pU4U22GYVjO+Lo2fNva3
YvwQ6LpdxRuGlyJHBt005XOGfODiJQWflXXRLuLclX5qMtqC/2aH0LtvKdjva0C5
eNnDDG+E0FXIR7NnMQF3UPU1fXqotxJvtLuvC7XerXLyN9MYK6/tMugGvZN/T0K6
hPvqtrcUQy6oK7m7Uog7NONmmjuA5Y9Ro80fmkGpbe1c2yYXgQm6Nc360V+F3nsM
X28GzfKZqgUvsgvDQXcMEKk5gmG7vAF7+4W8aea05JX/lqR+bosfLba2qAszypqO
R8VOiD6GWtnDFGdY3CdnRaJ/wEsG8bl7EG+0+SAagDPuoh2NAoojMyjRD9rAavUw
cuqg2MIhiY5C0KdvbQ4AuBZoE8gqwYshK+xV4ecmIFhTMOBtgZkapIG0UgRfiptk
AtjQaLdddpJsEnuiVC1NXE9pneit2IUXyL7Uoy8A/DBQWgBs+NJJUpHyDzlud5mh
2+R+Df/LgjI4uA7r2tuJqKq6pXG1V9d4BHjASdXywximwL5EgW/XJI/ZS8xng4GH
RiL4YJ4rouY5bzA+TpN0hAy7iSrWZyxoyKG0XGz7vwO14rJ7t6qZukVwYqAlyk0Q
QP6dYy/H/Cj7UNIgmvAMWcOe4+0uCSGoFRMKWMNXHtmQFTNjlve3vJJFpTLk3d0V
ixMNM2hdYSCeetDclqdYIKiB5UPpLUymPHRU29gyt3zkDA6tVm4SWPH7ssvURJ+B
fWcXTycYLTaq0LDyRSX9UhLmyewS9aKzgWY/39RGsjEI2M9L5Na9GVl/DpYOlcbc
rza49XlzDDqEukFyGLSic2soO/bPA/NsCG4CblKnBMhJzhSRdcbmjuCGpZZBwD1i
aL6pyua06qAxvUWyREItZQYQWqk2vPAk0xSUwFXtdBjs//mdRlQVA9/5vMuj4G1h
ry+lCjAV9Fmex5m/l2j/VJ0vSFF/dwaByNf+YV7zD31YazD1Gow2AgS+bFLKPwOX
/phme0FiuIXF8urysgt8Wi25sjx4y2V2lsKhulol8e43PmOcU0vqaYqlzg1fysIk
QWUj/ot1BPhxHkAiFY+Gz9jBAn1IkUBKrOC3ik9SeBUWODikbHj3YFogNHGSralk
a+dvf/cBMVPsSC3mgneT5uytJ6l7Bc6O/e0L0dwkCzYE00SzkTincmtEDUzhlfMC
/uZdHI4am7xSySNHzFSEmqONLRkkF2146BPZy50oOjCKo5ezZrTE9+eqreDXKYnS
aGwOY2X0/dJ18GHHI032OQYcScRStAnRGLqqI2nRdSBSnbatTJ2mcy1mMNoGqHQA
QtrpOFtAhs+rMkQnF2l9ymdEI8WBWmmNMb4RvoOZx3mKV8MyVMAmrNx0gsvZPPf5
ifaY2WelMxu3sqmALrHHbMG3U3138BmAf6wcS6hrxFJfyfifthALDQtdheFRUvJ4
ijWvbnliJriSdPuIKGA7uWgqxfx4E3FLmGoC5ldJSc6We2V6/5bIAIMGL2a6ttcL
bC2+w6bNV1WFTRyCaAxE0GNspeL1tKpUzqc6eXqXtv96qGXCLBYd0CXbYxsG5Hle
yPsZmotiV2Fkl+e5CFoL81x315FkakhpDJpF1M7W/ucIm4MoWl8pdjmPr1qz71NP
UGrXmphAK35PCLNR2P4XTyDpTvRgNaKAuscLgGD6EIeA0+qKg2yUqpUGfHV9USUp
SJ3WYG7oxxQ5DVF3sLgwa4irlgXwhZAJH5LYkQN2UJUri6GrEDBEQJrY+rbyyV5w
Zx7H6baG1JlHs7zZpuME+yPqd9d3GJG7jKO7MiobaKp+Z3fjDcH+bop8WuZASXfk
rcK4vXN8g76D8LZYslHjo4S7rtQQwxSpyS4cnBfXy1CeQdl/EXscp8TE+M7DQkn0
2tUZVP3r2ouNHejen3w5kwUFEcYK2V8HivaPIbtawrG00E0XkoDCs4XTkyB4Qwk7
CwbvtxoDU481udBtoX4puXfORBL64cNqD0R5y4AaV4egj3lIqSX89WVpjWNgEjNU
NCsKSBDIPg5jjliQsA3bs3Z+7yMQPHXuhpbqEcao7OxmkeS0/yaasOqP5L0Y0/Mr
GYYELAxY03BVu65MnmaRXxeim0dH30fNv2qjuaUzrZLvcyBZuP1nJ5OPZNnPruMy
oamTqVsWufJqpgy0A0Lb080p9gwscwgwJcI1zkXf26K8eX+x8vZg3ohnlgwB16Ke
lXf71QAlvs9TrVAcw27aMwkPzbfk71TKRBPI/MN7utDqASnlgAKp8oC8fdH5Dk/h
ezjUP+fpmWeMRSifqK8WtO1BKqMu/vYnGl78BYYH6NwOEEy9O+DUCgZ8w9XtbsRT
7TH9BYkmnHNaTTGlI6BilEddNP+7UHRF2QKBVDIi5mYtsdjVdnMatcx9J58yTpSz
IcUiKsH/MobmpF/z0EjCzsGu/fJ/gd6qH0dEPMx+WUDE3SUWgQACR5JZBQAFE8AQ
v1ldoGc7GVBTBr/vRVRlir/Dn/BY4pbDUgSDlnRqCFIYeBnXf03C0y4L9Z1fbU1V
REMbYDSx5MscPa/i7lAJLOSOP3wc9Uwp8ngnIWBgFikIFd+Uzk9HIMhwmJhjnwwi
g7pHz0fpN2c1J7WchUYEAROPsii2xnr0mEZwUKPLVGJgaaelhbk9nMZFJegclrYJ
ZHs2GC/tDZoiYHfIkhp3vl4SQTq3xY3SPBpxaZtAHjwQmaeoh1EuRvoclmtzWSoE
0tjO6+5zIZcuzWURoyjmK87aRmkw2IcjX2ewGZYvWWj8dP4mAfxnmfAgmVCLCa/K
9KlaS1bHetyuHRfAfvLPrqExVHg/W0GS3bpsJG1C6BH2gGy3TJ9S2nDfQODK0Lv0
cfgPUAaIo7oghjBNO+XlOGoJ51TqiTcNve3npl0ryhIamDBbwiVItqSPjfyt9OqF
iV5e0y4SDwf1J7K6vLFXeIip4RJtBEAMs4w8KQciJ/3wxI/emrmBMY+kYh/Zl6VE
xbRD5ThgTN3fhOnKZvZfHxF1szn2cYuxy6TPLKmWqU7Tuh65Oy8WSTLT/euYu8Of
dZeGf4ttfrtSGD6jQTu08q5dBfn47RnbOuC+3r+pDTpHhKcvLOkEbzUPDBAsEG3S
SD55mw8xt/4t/w+PENExc2akjgDZohaWXUh71xGflLZd/cf1gaWZjMhDkwOZ7jR9
KzmZ3Yd4oGS2NXc8OnWN+UVfu0mQdb0ERZyyl6YtG2aEKVuVEiAJ41pQrNUx4xiz
+GhPb24KobNbaD0rXDnSwubuCxisQl7N9hKVbEHUzk1CCUz4+mjDwpOqGJkdnWdY
3vB/jCZiYwnNVbn1y3jio/Hs4l900/W9nYDa/4/8KO5kPXNsN6+FCdvQe9ujk0pk
ZQSgWzHpo+3uYjW3JcjCNr9hjMsViqbS9fS18IvajzOAOZ2L5VjIyrI+c4SIaNou
8MIOGPldfF//1/cbTked2pVCapGFOKHSVnsgpF3LvMckQ/ugyyobnFiPrstnA5mP
YjtEdBTnHORnd6CXOrlm6jznnAuERVeW3OVH9xyIBNj7s3czZlXqH9UP+ctsnIt2
Nw2dOwmddhnFLi05ShZy/KyTyZ0i0uTsL3nxiMp853Me+iSYYnD4mYiW2kQ8/r07
ff+xkvyOmZVMnf3fL5KA+Ke+7uwp9RFdDnAbrORl/43u/5K6o40t0Yl0VbL2uGk7
PA+ZR5K5MRxnm/lQTXpgbPuBmKh8HPKflXNUg/FQ6/JLNm+D/AVNU3AvS4F5jRXj
O/IW+J72EXEtKYDDBgSwK2AyFhxsKO9kjXJARzmLsb6rbwNbHw3N+vS804vgy8r7
BtWct+dF21AFHHB4yuaiwbTYxNqTwetTGfcLYAF3eERpoDQysQcANhSxkBIlprHz
MdXdK6UANIQNw1TwjDRME++bz7nmiXotYxTSHxWKFo6GmAGQndpYklFVn6sUOoDv
wKF6uz+gWGXYY45fSx2RHvQy3PlMqBwigwWe+IfBQD/mxr5x4Y9FA9aL/+VV3/3r
ZD6h+xw3bLUGnxw0B6XRrYi8RANZ5FI79D3E3t+LuP8fmIvJtbj5MfMI/FHctsOy
wdC6XZPzIYIg9qfzEPapnRQVIYtHKVP218wzZMKpEdriEMYIs/ypOJT18NxuMoDl
X6nJskueITpOrg6qni+rNAyq8/Jk+nmmgqfLnucWabldVWg4wPczcLetQbACmHwK
sHc26k58dAKosNZs1pwuW2opOgEZRgeQmeO2dEb7sUgX1fitOUapa1sTKsMjHzZs
UaKSkKYpRv8xd7aGITHCMLFw1FCTiINP7TE90FRchprfwKJtc8iFR2U7lvUXADK/
b6US9Rtt4ZQ0rXe76IzwR42iyTw5QStlw4nvutR4xnT/zgiBOPQphmXR8/maQvrz
IU0qDwxIjHzCYk3PTyAKdmdJ2n8b4fKgwolXoCAMF4aE24OJVJHWF/ac+BnkP6+S
V2r8QyFp9cBHwOg0sBQzeBMN3rlLveUaqX0vWDedDs7nyxr+VceE2By0jCMwKYpH
kO86P+yf98Htvyrhv5kNHXD5odtwwIWJ8C+5hxzKNOKO+sb4hUTfzUbVG8Q1fzut
xUhhwr+V9Yqw//6E/Y8TpZY7b7gE0IrzyZa7FmWT38s8+YQ+O+v5YxnTZnZ5slyY
zqNXnl0wuqliGZufJnhnoC39csQEpqK9y0sF56+8g8W20lFUQqri2wGoUCE6sUYN
nE3k2rflV9HfNdILKJXIpLCFhel6pJ2EzaJisGjSi+ATVnOqktRm82aAQuSPT22T
GYFZV2w+X2AUNOFMm3MWYiSQAPRfMS8tbVpiUGJac2nELhLZaaCpiw2Zr03yitJj
SHUPXez3tJM1k4Z14tKs4nmJBjSvJti7LrQeuVlnP0qnI6SJq4rLxxHmV6QG4+sb
JOXN/GbRsyKnrcuaDJdnHKlxbreEqIahjijbcShbEn76kBZqi96qW8jdStZ/bOfF
3jL5ltrNgC73gs/g0Ws3agZk2Dx+WnU5/Hn0TZOJyW3cViLuXdQ0SSoSd3d7aaab
GOSadphPw92OzgTB7b2xFh7/tZAbUP/psQXoMHhuKkUo9YclVOPNJB2bkbjiAYqb
9PjpI6P/MatguaB7mRAyvulZNT6YnPIRI/y5dtE3MqA04JGRJQfxqgFqlxzzrqNq
KiYvZrdnEnxiPr142HOq0pDd6ZJxtnZZ8Sj1O29jfY/xmUarc7YDSyxIDFYkV/G5
V26x5R80vF+pMFcECHwFRD9W6VHiZ2Bp3gmIA55cw2hVbtdgdPMEdZ4EpD0sP4O+
KvExRkTPyyg0tvEynBaX/MrX9cfDpNkxN2eyrXUy1jC8VWCnpD+PQeu0V6mNn5FY
vJMe0T+Z9kIhebAKolJB8HVdYBcifYJUMatQn+Xz8eC8/IXUH7Zb585luHLbiHUO
Fq02X1j+EGWOjnCOe0nwWCslsQRV999LH7kQFKs4U3aOh5aG0tOuCF3J1Oezeg+O
8eOOEXnmtogkAqjcIQMfNQm5qbWWd7qydkzXbsEad4yYQvTeIg1XEakJIKZPY9d2
BY/dQxLcSF7QCR9NLmk2ZwLvXlRzZsP8xtlx5u44ppu/yGXP8ylQXAk1x+vDogGP
sZhye7ZI/B/sOydUfMW/sCKfKcSrGCZY4ZH50uQk9sCsRXtGM7SmytOhGu2F8J9v
Kp5AHS3h2Y8Cd7iL5v3HvSRhgECjlWpQKT81vnXRU3U4Zy7b3c1PALUNr+MEx3vi
7hx2PRzSnpIVPYlzZjXPUUqCYAs+Qnom5ByTbU4R7/klh/duTHz0/sO0/fO1XLWS
gCkkKYmQG7hCwdDEQJP0mNTxruIaiotIkQWRp61jx6Pioj3uND0i0VF1WfHuwhMZ
IQqiCKJBsBW06HYNGg7JEMwF0QEXyKoqbUjLEnETgWeWQVQ5CwRx82SCAMvrnyGQ
voJ+dUH+OhuOQlDTB72TZbLquzTAVhK/eP2QYuktU7hmN1sFNUbIUP4O6UGuWT5x
bpNQ6Tzih8YbHLxyfkmzgZr5TCAtucAZNr39c4+0qIBcf7UPZfX78RtOiq9LQZsa
iuG2Dak8aeCpzCyemjDh+X2vEMI4a5WNH3o7SI671oDDyNwII1J9ABxqldVT6+O6
bpTlBgpHUfVHUEAgYiLXqcZLXBcNAVIDCm3Inw9jNCmqFGLfZnrAsA4r4Sq5HBP4
JCrKrO0BQpFOYLCchFusNzF81Em9WCklGL1y0cCgNKi4H9Ghz0w0FUsxs6oMPYHA
g9vo69tPJTrVTh6We541q0wRLXpWXLCOYkUOMLBoZE/xHKDlR73KCpa0OL+8tRvA
w0xB9cHRlhRLjP4zKirN8olYZoYNkRXJjKsJ3CDh96aCOfPRUXWhytPElMFXBsls
clpT0MDSfgjQ0SKUaF0KLXF2GZCZsuRS6Ovi7KRpJ9LIKWDXT/A8etPcFRkjfTZD
6YPeCX8LbAoEzHxQ+3KZM426WSlTZhajsrmYxtF4zX3RhXxWagnh0i/dikoHkehg
mA9elLgSwIhIyNzMEg7c2dOurZbFWUAYe3SIUV3+e45MlJa/6HoeytIpPqFVfTmG
cJ+zRXUvJa1gf7ty63eylorSeXzYozoXGDFw54d80I5KWXflOp7URaCCLkgwafh4
A8uUOterdqBBoZ8tVyB006uJR4bZSPRevFZyMRa3HqRfOeMQpIuPWyB11wsijRjh
2ID1V0DvexF6sW5EOKoZ74LcmXEcOw7e+QFBL+2xo36AlrgUFPMnlcRwJgxiGdal
i9xgwz9hYXbV2JZ3QhIRyzZdAkrVp0H1RLNe/5X5NontaGwKXLRtIgM4xnfBTug9
RPWa/XrjzkMI0NPhaBGFV0yE6xDkEtsVu3HhpUsyBK91h4wu4S46gwloU4kwXXNy
2pWZW/vI5s9JMP8V9GW+Q1MjBWUDYIwTBJH5yDMu2bp/eF31RI5ui7ESFFa1vY2J
0Ud3q9XKQ0Ixhe6DAOgONjPY/ZWkArr5mITJetCpdgOeRjity+tbK8duRcjK86Fi
fd3ysuNk7yBLJIhuafNzBAa0PmPK8ysx0jXzDGMB0U0X3C7V5DRIQD4YpiIWqxLV
dshtmvLOYGmI4TkHe4Gp1GRrWW7qe3qH0WC/l/C7atJnEOtxjLLWa+kEnGj7KS5C
k1d8Y61UOu7ucYwdN7U2DBDktUjeymvUKp2W78S4UBfUA+R11G//vzBw2TGyXWrN
wwRKfCYa36/+0TlRZVtmctPgnqhjT8730wf/mUHTtniJ4Um9hHopWy+hirlre5Xm
RfXr83GE8asvp7vPr++Q951BvK6jZ3pkYhPv9kk9VVEeSavn07FnpQQAIEQdO15G
1hvBJVcot/1DCjQJfl99tIWLLfn73K97DSDCq+8Uyidu/satncX+TeuFW9SncaGb
mMNhmtOuGuqJLiVVeqkuSrBjDO3vUoAAgkZ6KVRZ1FBe06CKPGFwqQFo1fG5RzDi
MACZfQCR3xLVPlll8vCCQt0GmHb+Meh+UfRh3l7pTzBBBfMNcq/FRhYKF2N2HADZ
UYt8sJIgYSjqWHB8FJ+SQNWN/kUwstQwVkwfEsx1Yh+o4btLBI4u9BW9GweFwbW0
EmOxxd4S7SaOnxuVEvlqrGW77MJYTAmXYW9UWAERCaYzZHwwmdRSm9JaMle9t/Fx
OalicRD7bvZ9kThrzPaHJHmkiqx0T0lq6G9gzQ9wvi9p28t+98mhH68cx7dkWJBA
ARpw3QjkJU8M+ZEb0JIB6r3ohypxieDPnwhMhFLrjr9qY00zDzQSlD+6tmZlUkHj
/tYPDB6EFZuCTe+xYd+Ntwz7rR8qi7UzWnoQqc2dvFkCYg3bB4Kbf2VbLwaRPAS4
Itq2aozj0Ca37XpcNlx6x7zT7jsUXjnuZ0N9+HNbVByIUt5HA+l9papXpshFpVsr
VMuDyIr6kQDVtXEFyQtH0YqOkPrhNZyLr5Vqf7DVs4R3o3zhL/DhvzB1m/LJbSWj
mK2vAUmQaSJ5uW8NKczdZ9scpjt1QlL9+DZX3qhgZ3SIbJphn5t1QT8mhF4YgGXV
Im+unvGUGY4GMGZADYBZ2RR3pQYy8WqadOx9RPqFoWxOnMjGLUuJI0ruIrU86os9
Lgt2Q4OYZkirgICq3ESZTTQrbQq0VhCwjuCgE4blT1g7Ht5+WOBxVSCqZd2V6VRC
p4rLw/ZejQ6NBL4OfH/jnMpa2XWO5exbRPxiY5Om1KUOo0JZvUA4QOLkmSmxW8AN
NLjBE70ZXjauibUkJlaPWzOICUfaNnXOV5ne1hNI74P6Ns8iQ4JorZ+Fmnrntxf0
A18aXd4nvv1qu3gMB50sneIDQk0J6ZqAFT3OsKQfEv6TO0axj547kLIomebuNHBa
4GvJdCSqYXNjjy7jwMt9tRzDpsKdlT1xggpgL2IzknHou5LEL80a+PtYlG28fvol
zPEw9pZCEn/0Lgyy/RO3A6Ci+QklAz4EsEQdr2BxWdFW2MC8GQK8UMrFgPIBsAK1
s5PeWfWvphig0VJV+hPmR6iV+h94ofGnX8kqVa9QIfOwtNkEVvxQ13lbjd++8/7V
w+V7mAdoYv4MRa+OHa0pTG6iAXoesUx+/7MDl6rbXyJ3nQ+U+sQeGB4l0SWN8FPh
/hNGh17gWPHqQYvH2WXNDbeonnlLEUHgsIlXtQMF9fXiv27qurlOtUI9zIeHmOMI
7RqNBlI9Pmto7qzE9ALA22AdaNHi5LJPEyi4PDpYXcidR9GhYn7w9HS8g8yJJs6O
P0moL++AVQgW5lOTNrJtu1JOldsvP96uwbVmxdzT5eFdZiNARkyDnVvOKKKLpxD3
Ukec3/jfFyBiqmIg/1AcGqe4tf5kIW+ufonXtvKfYbzY8xgVW4eqrAD5iVb0qaec
yCprf8mSoiDcQrYz1DwxYRE6VxH7vcxuKunGoFAuP3NtE7H9hLq6vSsAqQ0QUrOO
CcnSnppzFl/6Jt56B+OdFs0FRjFit85jP8ESmZ4YtkEn2rKRGBHhLJuCixLS+Wo8
kFnR4zp4Lold41yMGomzhCX3bwJj7FE+vWhwz8+ZjTYnsWbcRCt1Z17liTQ6Y0GA
pCZky+mERvkJ8CFo75AxoDjK/uf6jWUSXVCsXK0s3aWaaEdWdnTJvVqyVl+V5I9q
ZyqOnBDN5RP96M/a2RP5ArEPWiDwOyHpTBIRUE5EhyNdwSbYYp+wFcufFCCMLx5f
DBLyGs44hf8JcJrJmmbrHETIO0iDGet6+C1PDp6bnzBTKYQi1218mFm8veAfOZ8Y
YrXYhOUVkaXBDtx3VkaqnU1ir5abmuT/O13tAI2+jwePWHyNJgyRBpVT+aXzZo6G
DdfY+3WDFdEqLd6eWMxFs7hVsUFGUfTqhtFYir4HYQZHAe38F4zTH8g3KAuHbRA9
RUGZcY3fcA1p7bBgWC6U+nBvB+LYfU/yb/rxnJ6iaKjawKK5QiJxNoaYf9BV4Y+n
3MLBQu1cWK+otcTkhUeY0cFRrb7mTQdM5iCIICiJLvZ/X5ifZWR6+EXryJqsmViR
Dc32L4terdQN3wA/0m/LeOk5AaWpLKjdC+s4w2SpLFCBRg531nfzFdOhwXO4Hn8I
wBThVnnXOj7/OcyTdQd/WQtnLXwrYDxJiNLVFB6hMYzhDo2CoKJiSqEoJJqe5xOc
rwNDBoN0ggIAoj/qtjryPjw2z9o+bgsDzVApY2uVgtGo3Eu4jpE/yNQMiqfpHrd1
ouclA/dYJC82QWZRbfwqdiWdAmmiJ7nfS7VZ/iqCIHI6egL0pRrlrZbRlPqkpJK3
ml18jYp2W7fhpI9n5DQaQnGqCFoP1r77EHb75bL6n+EbwyjfBJxR54trPIo9Zhfc
JQyAOigm1q/r9zjTpp2NSYselvsVMjsZCtIUq+/dnn9n3WeVKAWaycAyAzGHujmS
OneHhahkXZy6cdaDY1dssgc7LtxBzdzF1KHGzyoB3g6f1GQKvWJtNHcMNRS6dulB
WKBJdvR+RCH0JN7JeKxe3fYnmaGlkbx14lf3r9c3cK12RfQAKsgAM4R8ewiKBdSM
LCzUh8II8RQsjyuW2hLTooTek//8SuK1iRPmdGWumJp2To8lVIb6Vk0uQSaTWJdL
L+66f19/LEnYL3NF2CXo3e+m1dR6FFARAdXSHl8CpWzfPyjGdCuxy38+oar0aSJ2
na8ViluCedE2VOv+AEUKu9KDrMbHjhpJLp3vf95+3vg8OCzUZbmHKJMLfr7J7H2H
J7y+R4Ew2IMM4/2fjf0DrebCSgS5U/I5KafLXRwoqWUcTf7kSucz/n67+0LDX5Ws
ArMOtr0yMiDEDbBIfYbsS7HF0bofotytB1pNVmfI7ieX8qMoENczJFT6eDkP9dze
FX+vOzZn4n7t1UMBsDlGEV8Dm+GnsAulZhVHJ3hsezwVUMw0iIZfnrorzLOSHzla
TQQTShLxwhA99op3LrhaO2HDAY7fz/k2RgsqYmGj2MtqSeNq0g+IbndloClTlrRG
Q+Sn9PJjWDCUMhMuEKkjaA2EbdCHADDR5IVLobNA07gbnigt5n4uFcFXYjOyfrEm
BFXGoty8sD4UL0zG9YwkqKKXNb8712e0ta9URxK8ZPJeNjEJrzVzUD1FPn88g17g
G45qOcltUJX770Jbsey0VRWFtuM5bYAxipBYHM17Uqd4F+diDru3+fhUKEDrW9gW
MhCF27fB9ccQVRa2lybwbxLdoYPqZLSuIxagf6iwyo8bowf9PNiuTfLSLEas7suh
vNnHurZpDjDZ4Tr2vGcDQdeNX5XApL/lGj3QLnE/teA5cXBOXcVeiiYnw8AywbFd
osOqm4yuKzVpJkBa03z0pPF2xf6o+nMYhTo8J6YykOtsB6p00BgrjSaQXFBVtyHz
37QZ8DSFkkaGcKTfTwq1HlD/UJKSWPH1pc5ockAMb8jBWa5a0CtNIBmtwDgfi9oP
/tGkMsmP49Eps/fcdnIeIhmsMlxG9OgzsBvfYep7h2u+dzzwi/8J2dAKJA723F6M
KQwja6m9OI133p6K+qdVY0wAaCUggRluBjEk4SQH5D/SRNahl7qdgcez/gyLlflr
FE+q693VfWDdHZF0aLMU3gx9S8utJFupQjrrfrZh4O/Mnu5ClzsRo64HJni/IrYT
LSLDAj+Aq0AaD7dCVNMrx9Lrb7h+8wukFCHAvOwgH4BJDv6jhvl0cfLf4XfHQGpK
NcLpYShkFC8CtKViVoyVRriZo0Md60aW/DwA4oVm2GCokKc1dVVUsdCfHaeieq5g
T33YFBwU1xNF2X8xDUuZ1Zz31vZopXKf0S/kaxymWiVix61RdyYbSrYuXqxWS523
dkh2LEjc55Sv7GpZ25YFnXULf7smlXNMR2jGry39mqM2ifNdkbmiT1wJt5i8KjNX
HHm80xzu511Dc490RmTDuFaUfpcaGWoqKQSfchXEhID6LS/bVT/rjLy1hq0IZgxT
bwIRwRT+zRjJP7+rNWv0xUPjRImfKRc4eDxye0d83Q4GyqHuXV20S/q6YJQmENm8
d4hQ8Ub3TP4WOvB4QcTMdIz1pfNOf8xnCVuqdf1RTskZ7rYwlDFzjh1UwuPLEpgx
07M78LudBsJgC1MqxaoBYIYmFOsNo/c6xON5/ad5ot5J4EtCwiuvItNaAPnsL05s
o4/EaPgx8Kbn+hUSS9wZ6qkNpoZV+OR+p2M9qGXbAODFgETKz/YWEiBx2rgH7Mje
1Bvo0Btnj2ec/n2nYe2NRWcTBJcKX3sfRaNPAV1VDTVfyn5dERoeDmsJ7EzrivP7
13+ZYtIFeFLMLWPshcLFoYQXiUrraQxS4mb/o9AqlxNunRWdI0i9//roEXlXQC9j
0EE8IBiQqFJEBCU1XAfmDoCvWUi8keqtuG/jXbqYbmdfCkDFXuSwrQX1ujC8I7UB
h3gcVX28sExR1yEw9U2oLxZ31wf7RH7e6++/5svO8lpzCTYY/T6raQ05Me948QEp
UZzKtsly2H6sWgFnLhupmGO54RwVYOx7jl2R0lD/IvlJkF1ZGFzC8eeNvsaV9W0s
93qqdNaoPSUG06WrU7FKo/lyMr+ineqsvrm18OjyKw3elzQHtIv1CHIc/kzUkrH4
VOFd/Qh8cxl0MU3XBPc4KC50e9bjAxXubkBuvarfyLKLJyr9ZbufRT+g+SESVSxn
IeV0ZOP+fy/h6BoXai2FIKfrzeyKA2aIsgbQTkJdpI+o1F+H2utijK3u3mDzs4aW
fNV9tSHhSKfuOAdTwThw9jYur9n/mh1DK8hhyBMLgFspnZdEuD/Hm1tFnEjftFbK
m+HwEMvm8j8Y3h57+es7BCFQE8tM/Vj+FtrlTabJ73qnSc7oSL1NhrfWge/bn+QY
AFlchCYq5Qse9sqGg94p/LAl8BbLySdQB2YlFrMyKCYwy6PeFTpfwwwbbY12plgV
lABFMkrGq/vGk/QupPJAhKt6IkovdQZ7DdV5hTS7itJKbYw9cnGR1xF5R5Wi8qJC
CqUZTcpfV+bXk3vYVZx2d72Z9SGuo88/Y5V3ymV9P47HnK/9sj4+d4XuCX+HoamK
DUGVqT6JLWm3X2+YSQVLMZQvA5JlMum0/XyssgJxw1BcbPjSwaswtWhP3imc+YRz
97/FVA38UGfV1zB6JZ6WkzMK/4ADuD9JFKcVh1JKWFVFgtiGTFKZ3xI07wrFXo6V
gz8FQoLshv8T2k5xMMAQp/aRVgyf8LGajU44y6XaEzxnfiHWL1N0BEhl787txLSG
dA1z9CWsTkSTU0EzDXASL1x0gzGKZO2JrwvJq5GH6bogWdEOSxJwWJWgGo2r2aOm
eKCjJqqn5sXT5cHwoPmK5tAoVggtL7VlnWS9WsTwZd7K6PxAqcjR9uwMAv44BfW0
3Xu4rx5knEE88M70rGlbTHJ0tD5KyqEzMvhRObmpiJzhmTnz99LuS30WXrQiTp6h
2l8lGx6sHFpCTcUx+IY5Aracfbfzs6R9L/HDk1qXO8hW7hawTvV071L6xujJcA4X
Eh/JEpzsfZe6O86AmdBUSTK3J88pl1iygIvbcY0A7NqbrkMTjK/THvNy4mzRtvWR
0sD3UDaQoI0Lljl8FX3vH7/mG5U+/wCPaBjeiInCGADaKsWcoec67Ba2fMiO7k74
lX1HIn7hVhNMVZo6Xn81xRuE1Qkls8h4AUHw+eEF/VsXrRbmCuq25P6WZHhVX/4y
1ecH6Xx+datT/0Smcp9/tAE+H5Mq0nMBwEtT2jF7fGKLPUocspJOi0z74MkOyNHm
hwsBUJf/b/0cwWEhVEFOram3LSR98oPJwgJCz730jPcA1ZqcLucx6J3A8QzM4AMW
Gt33302i4mrmKy5ioQxmttQo/aHKS3oxEbdXwkGpI8vhMeboXgE4pPJA6pzGYAfc
mdbJZtX6d1qoTXxCLN7vDsQThcUFkQCfAtrq3oNl2vWB5MXGXRmBog2VExveMD1Q
J57N+14kU21RBvTzUNSMyhEzp5tr6iNYn07h0HScKIy3XDwBihPEHXFA6ZSegURf
TdWtQLTdauAFhRWtm6Ee+adufddIXkjV90eDQX2zW9UzTipsrsCBLr5EJqFMvzKn
AGLeL7CUxhxEyCoWsCJnfi9lQkxycw43dHEnOemKdhilOOOA0H04nyFUaUky6bUb
1/YNE7r+hGPfmTjKVA7jxAGAjqQHEMs9GXTYUo4n49erxDYnC19yKskmUh1dYQYB
ENBGocnP6dfmf//Go/HTEcCcfURDtuh6cjum019iiWD0ejtltGItb1YTbPkXVWCM
UaMjdijMWdMKPRAvKlizciRgL6FDkjLp8XUbqoX0BGOyIQBef17iafYTcDcPhX7Q
j/LWlVk5kjsEo+DjFgzbI2bcs0r7ki3OjqhIq+ZnAxrSbIAQkQoRWDSpWzT5iQNO
Z6Vq0PD9I076n4SutbmA48wjoaAPn1l4vMDdQ3/o0rFmCn/c7qNdLyKc6FHpYmlF
tV+zedf5h3ccr6bo/3Ayx9bMQikf66v8WSEB35VULIWklwTw8nLs1rGwP9dSopS6
+tL/Nb/BQAqh8R0C4LW21Lq3gN7vEraEB3oNBFDKS3KOIvYZed372CJDNuKgJVHF
On0RlCdGhhDF9pxs0aquvKUQn2coyEJeKJLJ28XemMQtIkJ6Wg0VB5VDY10RWbWc
XYBt1yPtcU+yRQPPGsz3TCGS5hXQicrVr/jI9KqJUHy3O3uqN3yOreEiKudPp/VB
nFCcH//VkoaK6dsrD+UKnEUgNEJx1Gd5EAj0EtlDqf8mH3NORT0yuzSaUjsJqD2i
IshPer4o7149d/CQwiiGV92j3iXCuVhrGDHSAajGwOePUZ/DgX+DyurYSjRfnOHE
8cpgb+SvplBx3qm4hDjFPkzE+p82GJV6kSphsnUVBuzISjEUnUTiWAvYS4dL3/Gy
OOal5pW0kX7zjdniLANqAIhZb2Qlpbx74uj1v3rU8oONfaZP7Rg35yh42vXHJhDY
ME0ULRCURegbHKbQepiWUDTe77ZYKlcVRvVoeVFRVXESCYxQB1xTLWzWaR4v+wb/
b2aFjDALd3ENLGJc0grICYSpluM1tO5+rD39wWKNo/J5+Pp6xN10E6Fsjds2oPF4
dhD2ubTINC8hjV/Icp4RyQVVfrDtat+T4SFQAYflDwEzkIEOep1GZpQq3gpNCo+S
oLKOr8WZ2fHxlId3q9WeEatRm1k40vxZttYtfnAY91R1joq2jgU9pali2z1BFl6h
ooCuowgIQ1AbdjtT1qxz9ra9/01Ho8Eh55cwrwX70i2z5w7eeQk+VMVFnKF8k830
RlcI0Wa2BTA/zByE7kq6hSVgRgjfj8qRzapObWhHcTXHxzZX0y34yZC0X31FXVLO
k5RXkNVajQFJltKfmiVq+jVzeBs1Rdmxm2eMprucHp1L9HclSxDBnVZSnkWH571F
U6SIER5TJ42xF1pWaC9EJBmMwDiDqwGH245CW1Ts5r8BmJAQtzK+dHgh+9rk7g7E
euV75WkKbgS1GvGiaYAjEJiPUXPFwzWHaX87k77GUbaysCgLOnRhJt88AJ2Kyz5g
0mcApeL0ue9u6nuBwGvg5AZY2GsPPFaU81QARi5w6tmUwsB5JYUczM9I8M6ZR4t7
e4ytvDUPmHWp+OBikmR/vsKirU+K/2hfALY2ih1W5/W2I9ZTAJvU50drbfKgvUDZ
rwT4w13LDiHJyt86yM5i7mj5zDePunfyKEarnIaObMVApaBJOqlX74Pygo36k30s
glYlsDDx4oYrj2aVS0wfBRGAwv+WSH9hUSGyWThl2QZzpJOu9uPTou3ohF82xddb
ecy+/QBSRhPUTV75JnXuzZLqg3+ro0UaXip12dIKSazu9VkY+GwHElLjdC8viDif
OdxDFG+AucTsMCkcQB6v7nbWdJxwNr/WkPSfwWgYVef+Jeycc1SLTZNnH52eXdII
mF1rhF0MkCXqekaxwicr9ajmHKL7xBDQXg3wH2D8a9j0Xm/Ok439VxaJA+cfrbPO
LgOnj2qmXC/RdyNsK7b3sF7kf8Bf6AfECVaY+Ex0b9rIDWUrP2R1zwJNIrbxDskX
jUfdvdtex4cMRk0Pmq+CTrXN9n+rENVW+QmZ0l7+QOlST+rJ7ObQpe13EcXG/3cw
JZHQCC7IudMA6AulN0DmzwU79PVNV6xcnnUgF5HKEDbvdu0I7efSZlhlS8+ah9yg
pIbJit4zN1cJIZ+wj6wzoKi6XCEyCMO8ALOf14dB710CTHHKaC0+gkYwcDSJS0K6
P8+GZ2C9N7Wu2NdYhW2dffGH0CcKm5GNBCdY/egZvrD2W1TnvbCvVj2BhevBnwxl
d1D5DXHnDyP6gS1wXnujSeqVAHF9VGZV2jap9L+YeQRORN2fFn55qNM1QZUlFcaY
aSF3fxoNEk6fo5WtxddJo9htNMOWapFRygvA23KIJIlGtIZMJT/VMffIOB8pWA0E
dix1kKcucAqSvCfAhPe7s3WSxVJ5LUin1Xzz4LwmoQwM3XS2MRznOil6WDmZIfTu
sj/Vzlzp6+VgD2xTxFbiI+y56LGCybAn1Dg4NterLu7KBh6O8uhjNtOU/r68dSgX
mPhYcW7ynMNzf1g6xgXEVXe8/y+YzrldFbHdNR5Pey9vO9F1qKxpg+1PJWG+uses
R8jPTLWnocv4YrdHW8uYP8KHexuK9z2KP1PTB9kcNp9idYVsLEI7SMZMYMUZ0T0D
YKKZxLkLzTO9rqheQIaXN881yf/wLKDcOb9SJcCAbfVr/pb+e8fNE1l/K6rqhwlP
stGWNCkhPgJLEvHqa5IWvPz5CRLT9UW4VQDVclx8Y1/V82GP582X5Sh07pqGY2WW
meNsSIoew+iPRMFsSiW2mb4Sa4+81EjMw82GoHZgViTn8Af15X9Pgb+juzuvmG/G
dUjQ+S+VpkpP5F4Wsk9bpvXQdx94UzRppHmYvezFib64AqeRF82AJxJ+6DNeNWbf
+UEmqA37Ogo/eUCJGLI6KjvGMATPeraTlqLZh/E/+pYMx3GLmZgPRip0YcJK68Uo
r8SjS6CfLrtzJcp31akVcBWRbOeyRsUM1mrgwFjWRtkjxNKFnXdsIEPBsnMSct1+
QZOH9tjFWVz8hlVdtoK4gt2DQA17mhvqU0lVKOyh42Td7nVrbPPMS2M/p6b+h1E9
5CItHqtBstwzt3bv5rfZcpSuHFGJDnnDhP43OU1BWiNbkWPyu/A7nBR5IxZ8RYsE
iWH8PGllP2M/pSi4MnpdtpENMuOmweyIek5AcymMICAEWiXCY8m+S6loYbFY9kGx
nWzq7bKcRI5m9DL8l2WE8SBxRsOzPJVYNyg3a72mlhwtvfhiM/1vbvVNHTFhZz8N
e9+YE8MO+cdSo16QVsGiC0JT+DIqfoBKoNRbJ8QlW4uRAAh5K8deo26EV9IvpEuf
4E1M7MHBYKx6jtsJoPP0HqBB7mh5v6DWszCX78/oj98D2MmazpJlcP5oHH4o8Tl/
aRWL11T2IhzLR1ovWUWP0KwD35ph/1yRFz2Wj+AJidMIHoGQx5qXzLp4Md/MBYPU
xCc2KgvtrdyuXOQ9+MExJrQbRZECC9DpE+M4xGlA3YkdXvdpqUC9btwtWAYaq1ht
XK+5xTOdKf4CmCHrIdN/BmIEqizjgSpoCt+leMurpCOamxlBNheWUYwF7LFGWKAJ
85wWf4m+4AgfnaWpNRiZTBsTYmX3/e6B/S3w5gDIFd9cbpYjd4U81XefECdRcRUH
ofNA0Aq6bnV5vxeXMkzEcLPTy21WIed+k0eLlIfPuaZhTTGDs0nGhUI7w8/WchTf
kIU96Ow6LZM2ChftKHCVd+JO9VxPQhSqMQtaq9p8k2WWM90y7eeJF3A98Xyu2yxr
d8cITjwZdNEkzcap3TWk0vIrloQW17rWbKJWOBRNHPbAYlcu5OSjpeaeDlqcke1P
UdTeaZMiEDox0a+ysDCpyXdrDhPoKwYSPG/NjyOcYxXrDfKQeDGiyed6TODpWYjH
dS9mrKoOdq1B+biIKx0C4chNFE0Vpsrbx1w8n26/UcfO+kDH55A8EBgZoDgoPfKn
wxSe75jkiypX4w6xqA+ymxfrLBPaNeG1NoQAGtyzLfuHyfG1QWuX/tF6ZQjSBdKJ
d38L3vgdbG06Klf7JVxhz5bhGxohtoBmkmZSnsJ4Uluw3zFZZHTvPCOV6KFcUroE
t9C6ebMLd067ytwxn60nd97MVkAMfCkcDjJuZr/oX5HdOZTfRVLt3h/Ncpr8V6pO
WZu2I5EL/w/YJ5Er/F0FQt5++m+ib+5vKzIPZO9Dw5tJ0silleYgwAaKJtJu3c1Q
7keb2tZFUTlqIg6johip9QZklaXLjMIWTlFGO2fOAMkSX2lYwY8NHavPkWJ9pnyu
y/0dsyFhVxu8LbzBG9vJBRT2dJuOa0rg3Yn8SS+ZrcFXsNvLKEnjh4jOcIRuw9JE
6TkSmcpFTf8buzJh0DCOWu6De5CtMeWJkotG0ebXu5RuvqrGyMKTw98JmOajwiYe
igwrBkwLDHhkvsyIPU/VdfI+CneI2It8o18IhoDrfzXESymA4nHnYNjJti+Ia10L
7ZOSehFYS0YhhYD/Lz2N+YQUlTXXWbD7a/Q5DmgxcSmOTDz71eXxpvXFAbGnXbkV
YPjujS4u1XmqbXM7qbXG52fO96R1kDbXoRZvziDVC7RXBH3MqKDyWUCMylpGB8gd
MUQYfcbZuVlf8XWq9Zj9zPEqRRUJ3V2ZasQimaUk0iEi3bkqn5PjXbMco+Vv/Lsv
LYxEMY8fBZlHZRSO15IEWnHMbSYHFjYr+xbSpJPCZsi4royo0Lulxqi6vmV6duqj
fgXzH0tqQMKULRY3ZdIKtATXOBuxrZiRgPUmPkz4nEZb2VRO+pKCn6dboiu1xCLP
Kv8YN6yGh6AMrl2KSkjRMnOa+hlvGuyUGMRKP0a01wLvs7QUrGiHQ2pMi0cj4ICF
9QGK8KOuWN4huuNsPceMKxCjpjiuSw8AB9ace0QQWDdKxzCYJ/SrAJu5MW9Jcx4O
IeNOkzciTrVvqBr4yU6Flqx+FXjsHZjM96gxW52Ht6BR7zclDstI0gCh54IA0/j9
WZx9qIK2gfwWYXt2sL4L81ymaDnZPKKwxN3L7qR2fOoOnBIH1wVnO1ozgxIoGXx0
o5xjTEyfZErisNnq2Um/tf6LcInbNWOJV7+tkYqgGfM08SmiAUaLHBhrTbYEo7EI
qZ7oBO01ryQIDZnrOugFZJWa3dEDbQnBMOw9cPLzUjYnd8Wc5/D4b0YOWf/Q6tpJ
dQTde486i04K9hBNx0wQW9iBW+D2dEE+ZGviautEJEfneGaQtjMUl8tb2X1nSAVR
COsNC5CBfEG5Fuj39DCWF7+MuIJTxFyDnwJPgKiyxRyLO/ewawONfnR0RHFkN2cW
LFetqDLH+DURZIBBI+DpT2d/k8jbTk9kchrGLM2yk9qxLHssNyuIDf2vTGpnCKyr
BBQedGN7WB7xVr/4m1wYov2xjlf95rUJBMkcsRK1ivwlFCHx7SEN2gFPlg4zxb2X
C6ntIkj8yqdnKYlif2DJI/YBG5+7IY6cpFy0jz+QbvlCghkMc5I2zu/4xHcuj70k
aRKMwtRVkJ8WwOqwKKIb15AFixpecp82hL/9RpNZXLarXajJWzSmfEj84k+C0Vg8
zZj0EQv2ZZ83/alI5I+cMIaq0caWIB0nDBh1YRQ09LQK0bkrNkJ4RNQAVbZy6uPd
9zB8N96IGIsQJ0ClT8jKJG1uvKTbmaSWt9OjkqChOokFduDgYDieE78Reu0XWrGB
G9y/AvMgK7ydm+GT7xQskD6Pn00fp88zNdtJm62Rro35oFD9WwGTWURpyynJQN++
GzPtcI4RInJJxv42AwFD9S7qLTugbXRhPOqTqiPrVQf92Aqd0wqDfdyVpsIqvDpt
y2h2p2REtCpYazCLfKpQ+jukyZWivIRhnI+4QzQ1pe0Zx5V35tfIH0e642t8+7Cq
djgv7zHDnwsp4+fKTIMlXtB9vJwYpvDFPBaj5FTAayK+SjAFCuS0v3sf5VRrZTe0
nwQf9pcTcwDW82lsn/rjgclZmXgaA74zwMuFB7kXx/v+QlTveXfc6wRqWHlbW0Di
oi2M0qcj6EqWxhkkoO3LHGeWs0Fictj/iwxApMkB+dxRWSosZTYVo5qR22W3Ab0k
7FyQhhkShPpX0ABbN1INsiG4B/h6BceJgEbynIjyLO4ETtaPbpSQJERrwPIM/85A
pcSoBEPOzUnKYEZHi46dsJ/LfvAFiTbBdV5C4qAJKTjuy6DmRSPczAYgp6srAzFk
lUamknyN7aXya7aqpATWhIxImpOAtrjjDVdX2pDtcpdy0RpQCtZTmj95GThFK6zw
5Y6sEiKWSC6XkKAJ6aegpfy9Wv1Lmm0F+3UzbEyV0sj5xYSG0fOJkOKyQchL5ZRL
59Ihu+LI6hWlZv3TOuqD4c15pVkPc6UFUhyK8VkTzDLdTnkYFLVGh41lDwI8VAe+
VCEE8giPzFaNrI9G3Lw3/XhiWKYA2/3twiGfKmhlfHutuuTc36po3lEMY6xHQ/Ty
GRVBJGvhRGfHq4CSLqvWWpFP9o2x696mOgfmxMfbZVAEGudPO9LKj/F5uRdfXNM2
PenVKz/kspEQcbKxErGnUbWaXBwUGSPFYByex4E9iBgG/ZtoN1b2F1najCJPRZ2I
durwv/tqQCjJVkINfwHKDolZSja7JOfm/ojs7Eo4dFXxu/qGONZEGcyQcjw09YtW
2lWXuzdG7NSP6vGRUfdoLOs3GOzJ677tgrI/r4yYxKKKcPahKKoa1zVXfvlwwu7S
fZOpr2IRJer+StcClgIa4Paxx/qa3Xm0t88nG5aLrXpToTl8Ohcly0T91qzFhNnr
vAgsMozGepjtIkHjscHh/b3DyaWFqKt6rRBTL3XTjJya/eXdhaCtl8Vtd+Vvlmtj
ubFJ0BHSnM/iEuyNm3w5QTArkefEsZlAdtEZ+yLwr1Hh39f8JzfUCkxfMNssmFSg
57UvugWXToAKs3AfpfQ+4BJbHZhGlQvsesB+9d+KahjRrO+KYXPTEeEeslio4Hhf
ixW0FVoAhTE4X6ZnuOnESntX2DUh65bj8gViHklWUWFuSLGVdF23uz0TGjhS4gzt
GKa7SQT0ORKbIogcpOK3WT0n+A7LRB5D3qS+q/+GzLwzoENJMzT/kvBhiKW/4YaC
YWUIelH3h97Yj4IvPARmUJPEKE6lnZ5RmB+GXTl5q75hCH75R30RlJ5uxc9YI/7f
LqS1OA0vzvneKt7Mfql0IRDMXjXcLkI6BJje4E6gPvJYlmXlEloaMLRjQ7701z42
HzdaAMZ2upOyKpHutHJGrI8kSiWJlvgQdj+GahplhZNxBFR4Tx17dXhWKzZoTGJY
C0ZmxHgMB91+Lqt+z6LD7WNKuONQbsbeeHDUjfONHowuHlFk+yj9mPqWbQylY9b6
gkY1s2Q5Smky0UoA/g1qHG2mTueLHkCe30mKtoCxWRE41RDGJ5qOPWB4wxNohI1W
N2+FpxfQvZgDRfVTvVvOOprUPFP5Gc8/QpbV9holTtPjM63M9UDCIWsWT3OVFwee
W3ThS2bevqGbtkNOsyE8Ij1doofMl6noajTyToMYgDB9wbW3C3xhJ/zV5wfB6eoy
xLdRD0FnK73GCaIaxx2uD90+V6ghBJ7M1gze+8ce8razFdFRPi7oKUhfKU8DW9JD
QbWXFNlhiNMUdkZF/L7A+7LoEeU/013ja2gZyd0G0ifhuSFkly/ZRnkk2uRl0KRk
q5XQmoEFdkLuoy1GI+HFGN458lMRNJBfposIDKXHx6gyxaQPzGQYbq7u2mMlmvuV
KYQ0Sz00hDnSO/Z8HgNeCXH7O1DADsktxdjLxx46XZDG7h2VPMIsbrOQlCHnYwmH
O4zhTOZMqF70kvbnBvMTyITajl+plABtny3pWF7K1kmynkYvgTGdFlczuW8iJSyd
FRzzSmVwvtkEvciPdn7ckvYa+zIXLSB2L7Gbi8j2/NWoU9CiLXOUEaaDnVXtk2dc
YR99mkbkixd0GSmV7wqCPZ+tjIVN4tlj4E+Af7TV6GEEyG/t3VtyIYlSMy3jjI6Y
p0sw2z/KpIKoByFR91fdojaj2q5s0NnpXAjsw+L4jRm2nHIg7vZRrZy+h9MAVIWQ
2KxSzuT27fZbzLFRZP5pNPjb5t1KJ7E6nkV2R4LOKXXy2iVaQAuXi2rmGsjeSgXd
1ETxbifKRNf3otTgubxPQyn82/I1MCgkj9QS3BRUe8L6TiQn9xzpWGO9KhDRE9Mt
8aCbzqO5qhK1fghqnA+0HYVgSEjD/S1QfnGiD2qWQUg8KAUmy9ROEVgezXZI8ZYB
/dfx+n8ZbQ8UHRFX8KEd7tnJT5z2uENAn1AXQNsU6GKMXBzU7KR6s6BgaOMFROxc
XmVIud6veqgJdYOag01K6lX2eaX29NDIAU0Vmpf1JpLrHr5NYHkZlnhY/tyDmjoq
PM371ioKU48o56h6gR4uqZeXpo4nbiTskx+oiHxfgm1UWjjCTC/7+sWMF91OyjKp
Ra+GeBzZNeBqq4D4vyM5JW7b+ZcuVyvqiTKDrY4L8B6vWorUWatTKXAWGJMUj7lY
R5WYdsCBDauCQ8P5H/wFhV8NL2kzpvbqosIKkM9B0Lkn7/iz5AVZSDFVUtz6/waT
UItQU6oSHZTsIzH5LkZ8CuCUZPLObX4LBYWtqdd9IRhRgBPjD/20u6XgOEPzKVz7
klWLSeOvbxmOTIakeelim/1r6Mhj2gi+4EGT8WKy/hSD2mRFmsEWlLboUanuQAbc
2nULyk69rjgG3I1APp1THT6CYT3mrv3iO7AN149d3WVHIouStJsEON/6w8u1iyIV
UmtCdGpLMLV4EOpAjffwNjay8VN0ZjLj1ici6sEVCjcKZyGbcO5LoviFafM1zCad
zzxfFggo3Tx9gCtNogBBOGR1z75zOQYlng4xKJ79E5Uzf3Aq9EwfUlhJlGyPxMNf
yikznNoNIyqaSEPFdk/PuxuQTb2Iav9XMpxR0qQGyCw3nByJkfr+oIbUrN+nNIln
NZDovUHM6mM+k3IcpOeoyh+4xDQDiZeQ+vixgu8sZ6Xgg8az6RWHFiPwJkw0BAzI
9abSzIKrUskDJuXeBBpQpJBluawewS1SrmkMd8ZJ4FnjmNl75ZUYprImqdNKEoHr
qDOo/nOj7oBqht0dHnR43eJTyYkqRgoygdkwY1GXDOSYK89W3Hfs8gMcNMOfDPv9
Mi68oS0lcKE3zDR5XsFQspsY1hOcVvbN/D98L/hNZlYOzJhETkcjsta6Q7MpjYHv
5sY2EDbXme4XuEJYNDbPVG3GOE2sRl3M/wIhAnvGbgEl4j+Pp4Ut8OmfgDRSYXiM
rn1RNULWsoIIwgWa1m73asypof61qgvWSLX0446xyfCWgLU09ymyN+XzYLxkdNjs
QpqdycJDxmCsvu4b27aaPaL9IfYeKdBs5/TJsuOryc5mLKp8ZVm+K/+IXBF6mUCo
3dYSUdCYXXfvje6AYZyaJ7saTfQ2TkUPnWyfm/imc1p6A9yK3h8JzHjXYYoqu42T
PANDxV9Fm8OfynA7o9SVvuQj6q31YMPSThsvnbIJo7WsE/iJ0DC9Vjc3pChcQKja
K7VLNIGNeks065xPQCCsYQPAW31q32LKl7jwKrOzTYLYM8RiXQp2m7uJIxkLYwQ9
kdmaqGSqSt16lsnMOVSpJvwX84PEa2OTT+gdyS65uJE2Gv2AsbBzGTwKt2pspsiW
6rXmx1j4cxNh/intmZjgvnnnISVzBT+pdAuCUSfB5JHyu4s0FS0UyC9cfNV3XwxP
prx1xsOVAu5EfScTF27OHVvKXohPNE145Fi4bF/a6em+Mnu2m7P9lbEON1GZZSQd
O1S4SQsah64gpX1wWmPg8c5OvUOXdQP6nfQv+bwZsZnLNW46UsHp4YQNhcQfevbU
PAg0NHr2aNGfh55Lpx88AJbvlQU9zMQzGYon5Gki8eN+WR97u7CUGO4Gpt0ztuhV
zVf1a+gQy7Aklo5ikuuohyuIbSqHViug2nEgl0aYMSbfqNRQRbKKziFzy2d+pcVF
9TeUkg69vKwUmcMcixSudHwDZD7i13N+Vm2vzFOhRTOE5wkQd9hGAuWhPzzJGzk6
RGqpqUt0c3mPSTYwCvPKsa5SxQK47Xl6o52yaitZdsqCWD7CvKq9TBnP2VMcp1dd
YpMTYfutQQZiTZOq6tWq4OYfqj8773h/iLV/MMkWUdYDVRU9CYx9kUETSERtjaQ+
w7DB4I9PNiZvI1oA5GFGpneL8ZkIhHYClDuAd0+8G3BZBJ2pfybzKLDxrET96UzV
F32d2CDXRWpSk4LodKX5LwLn6OS0ua5H72tJd1E2s8gUMMvOtDQoMPac26wTaDDB
3tZBc6jwiWkIKlDtj3QfGTvOI4CyxZQbxJU341tSI7Amyz4hZ/eICz+kx2LIPut2
0RAZdLa0AI8OFEn0NZ3c7uktCnWmxvxABXpj4ggtZre0GVAbJSk1U9U/vyg3Uoim
842AGuBFBh8o4eekEBb9pWKd8nrIujdmh6MABhLzclVIR/sWAGR65ozcj1/y4+5F
MIS5hOMZjGj1DJ9Dh03cg1tmOoDxGbnvF3YA5crz2d0g43LXTy/SVmiAVuQH7xpq
0VZ5YgCZSz+6W2jv9FY/W7k9UiuErxDKv9s9Ar47DY66tz0+MmEPcMfC+DqjZInz
JG/juomEr02MEW+OQSEV8CfRKFDyUTsYZqDaoYpv1TGuf8m3gNxmugRBXmVWwTlD
VibjqrZE+3xSvPqi14SRB47R035AxxDqVy+2fZ4k7Nw75JLoH/GQmdRKk+ZDaTo8
H2HNtdo+EYSKIdJ2Vq8Chqo4bsKabqTmJ36S+IlpFlMcz3K57HXtgEispPMCtkDE
TWU/MsMTFAub7Ifhhi7Gb0y42V/6NMeW+AWQlvwmY5thj6fovR/q+aauDu7q+lBh
dISdx2phS14a9KSpuK3goyPinROpzUqyqvmtb0RcDhd6fSbpcL5n+8+BjRoCdWkJ
pIsfMrpHwSSQvfWOmQcgUUeKTlBfdXXsOU0lHEpTiRy5q7X4aWzlfpis69YHiLrP
wTxppQO03wBtNHTIz9OsLNjCnE3I5VNmEl/CTN4t/vV0nTU5Xk19VRZUSA631Mqi
62/hPNCqO641QTJvfUrOUrM7zBMCpoCen7PnM9F024BXq+qr5sIuiyVdevJKCYpj
6y0SRLZQSuFr4n4mzERkwuVPGVoduYHReZD+2jOvax2l6XAgp/OZTTXLfjHWnovI
Pbd/HzcNxYqNDmEdgO8v7WEHyv5iAUgE58wLMq6qFK1Q0OShPa201uOUCNgWdHH0
MBwBgFTSHgmF7fqYJOO0CWHqldKq1Nc+XgMrJIgorg60ja0IIFP89CSD6/rJDDrg
DFlPyGh5DljuWM1/U2adD/wR9178Pknj7s4qTsOGrXGWTP1/iIKHiazPebLN44rj
JZ06hTvssXpadzvN/G2jXMvWZk67bYeuR4oEzqy+Cj8lPrzxiNuhyqCWuXx2xYfB
rPdig4eHVrdOjMoqPIG/mIm8yal9Xy+lT4+G5XY/H94Iva/6Y2Dl7t8kHfSy4why
w1xuozuGugGTAU1W5YzA/qGOEmNR8SVEcUrDniGEG8KqeBChDHaW/53ZeZqXP56/
Ydh0X1k+ge4N3nME+gCVnVc0O1VNPd9fjFALOth7UNozFjMZwFMXgiWjkgzwf1hX
d+H469hHhZNFGvXqXXmkJcOPpsJCwdiit+nGdzMZZqpNQLRJs6LJ5KbNgFp3WA3+
PimUsviCzpI2UtAhNqkTUgqH/Cq8CtU3joa8WK6QwwbhGGM4230CwrS+0RCf8NGM
GFWuHKXBYW3UBQGt2Wh6K0hwRLil5m7eiwpHg5co79Zbo7ramUeaBkDnrFOgmP9Z
1dH1LDk1i0kT2msfB0eSeNfkPdSYrTsdHz3ygvt+4+pNcegDS0+ZVBxleZtP7t8a
OMLU6IqtxzzssvcJhG1zenR3oaCAXYXSpZEQZNM4TbG5IdQyJ36Wwr0HgNwK1DA3
Q4RVY8qWeSwYnP6bsxY5yh/z52l/C03nCLlsulC+rzhBQVqlzpkT2wv3IywoRXvO
apgSdMGl3d3yFq1a78EZUzPHtKuq6YHgJYQMi5okeHiZSqnvOL4o9+uOa/g0Q/Qv
xrsf3p3ZIKbaRUCujI69hQiec93TPFvoUA8dR5litEdOmtuqWXX0LzfBk0GN4+5J
y7wSaike8FdFvPgQWbzGc6eKXpTar3/EtsGSh+XinIYaddwPMvJjd/5tJmuVNhZG
uvy/DKUa1pkDAj4eBNVuXOvdv1Z7zuo27Yx3zH/zXidLaiqfqEdsD/bflWJXNh4j
VA190w9Pl8mRml2iUj1vr/3ZNjW5pqzINNfDeYyC+hMU6RoN5tC3K1W2hBqLpu2g
6MdJNvWo88JIoJMcEHngPHnQgY1uG9l36EvPgaVsVmBpEvSTWqxURO+deWTDpMKF
LjsDE+TyfYRFulKLYaAB6Up05Va6tM0fHaZjvtFnc+jtD+GeHj7xsjw7liDtNHoq
D3lrJo27wfkIRWaJoZO1jMCzlsgcpNgXsyx7tTMFvofCy7kl4ESaxEW4Tw+Dcd4x
6DZkInzZKvTjh3m/SmWK7Mvu8bHZdNY4GCqAfa83LhoTNk0Wjrhwv90OerVGY4Wa
UnbBQD+VB2OuD0Vdj12RWVdoqEDuH44InGKhsE8qgybq4JZ+2VBwNxx6R1d8nMVp
rIT7f4/2MM66KMd05bIVeXjITstZ5T63Z7GvKRAbsBdHTu2fONP2hsleYeioS3sh
6rJzWvK6OW+0ITGnp61iYQMiCKx8Oh30YNatrVLPuDP81IaF2KQ+QCq4+UwjIncb
jvR5slvoAa8Q7hM1DpjYRMtZ7BLsBDf/hRn6GxQu/7qNRCveHjKlCdmaAqMnYlUk
5E6+oJmKszjAIWJHjde+xhQU2+w7+wM/cC/lVrkUOQksPIWQIXvHKbD0UseHL/4J
q2p4KncO03ywWbEBsu04qqLT5sLRi0MyLt8WC3aSWynarErd8vb3fdW5KWYqv1ws
jAt5UGc+dSQQS+kVpyPwTYcE0LJlHUYdbdr5jayO9ZVcEhkGAx/StyqzpELqEqmM
BJ6j742BIL1g18x827waLVVoA7V5Vrp9IxJeXTllr6AoXbD3m1LXYmTCJTXCtOtg
WQ+2IzGo52Iay6fxWbOz9u+kvqVSpQ2n1yDzAxoA41w4K2LX8vOQYoQyMUZEAzTi
lNIZv5BNuyMQX5q1AmH5PSut0LXIxvZMw+5EvMzCxRvzzJwNqmyfkQkElHh63abl
c9oX+3C66Tm/icavWjwNHCOrryHADvI8VnYztDsl3TEKhsIdpCkjqkGmOVrgr8kn
h1xXRouGQdZTeoYDQ7ISleZYrg0PbmuNLZ+QZXeh+Wq+H/FaWWqjtjRtVVCQGs6e
D6yYwUgfXZZfE1ZKR8iQWLK/Vqgym4av3h1Qc8aim+moiYaXBg9Gt9IszYHtYLLv
kIeNxRB5uBFkeO6ZJvtgYFu5ydKb0KauEQoddmPAElQG9Nl7IxYAhfm0HtxV5EBi
+tv7zDTV3Mos5mvAr7I58DzslbTLSNQ+lfauC7GY62fBRcbZ45yX9lO2FLPRyA4t
HVqb1pAOpyculrGHZsTSCMbyY0LfxlH7GgzFmhFLgp1OhKBrjBD7aDvwI712YdIT
8xQNRzBxF/GWoyf65xLwBFoNajyPjLVwgkrhtMS/kUbOC9ecus1HdaWH9mQXXyTD
KYUYVjFbH7oLRv7qT3Yzim6NpRsFDZ4qt2bhO1m3FKssF97laVnRdgpDUrCsN0Q4
kANZNp2Q3/sed9ZlYRHy7i4qtkYqs6NwFeQakS2hHotinFZOiqARlipakAyNwqw0
o4B+5JpvVGOmedyvewJmSxOFwNtHxk27SLqhZU6wkx68+sBx/w4TmwicVlJc4uuI
tJu8bpHKLkOKs/n5etH7JaHu8NcXsZYKPEPRHRdwj9z3wJM2hDXMVIlueMFOTKZE
dLJ0ZzatgmxD/FYBztpBBovVonvQZ9VNFNZNy11RTvW383RRWRbCOzfUA+/NRHSy
U3kslHBbJD+8c92pgTpIr02Bgu8OGEvrrzWJ93qTW1aqbZtvsjTsEY/RJKVM17/m
pzs05yk3ScyqpBLtoqTN0NfyE3fHlHhidSBRR8PWzm2JqZ7pJRj4InA93WE9nLUH
274DyE8YNT1JCxOR244PhGcG+usSn5v75t6d0rd3zACqtVWXz2JKmjZ9AVl6HEm2
o30DGHuOw0s0vHoEg+QSaVA6jp+Uc0iFCzvyPPtGsHcxZ1CG9pgQkrHep4tWFU7T
HwxMbeDaghCK8hJEh3HGLkmUBKjlyIODftIHcLvPNZzZJ5eCP30UzyJmUdL2ZBnq
X8OCtYw/pExGe2lLu3avcUeb3YQTYlmxyJAw3IGVTyl7+mga8MVW8/YasTnKkRly
zgupqz57OqaEGXeugNBY6HMLivKCT00RbWAs7aDkSHbWn0aRHPFo5zn2JaA9pEYJ
dGyPaX+ePTrgPbXJSiOnm40eSghXs188/zuJC8pE1XWxb7kB7iI0ECLAxpgKbZZS
3rDvX4ybIWcmZFQDe5Tzm5CDHGERhihbLbDVn436XfsQ/IlfB9HHNBhhGAbRySk+
ZMqvx2L9895nO9Dffa+O8YCwGPV4k98t5SlVA06iklUBnELLxAf7qvlnQtqxF0Sc
nfwluEzqmlQY79ChuMjrCwUv5fLkdRbdCZ5TuJvMsVv5pUhmLe4wpZbbUO4ZLQJ9
ZVPENeD7EXqwL0E/oEW5cO4f4Kc4Ew9t3/5TWWuibR8CLYbl9+f537F1llo7/q75
a09XJ9xKBa6AjQGa2FT8W6PHK0H4asaM+VZsC4Sk2doA48LBkxZfpjJhBC48it7D
XKH2AcIoU0wy7Iisd3g6ZDDz+moCjNqthaDcxR10FvGycEIKgRiUAD5q0td8cJ5X
JYGGT+txhftfclj2pief6k+qjcSQocSxwDEfugr/Pu82IMA8gSm8ntOfuua+XwaZ
LjLt9p4I9PRbFlV4tLOmOPtUg0tyMg6BnxWI9jelWkfSVpovuiaESauRdhu9phf0
NuqijwzISyeomFzK6KH/gn2yO33n3wCRIRuej4hp1HuhCv896jqO0TAfN4roK6kp
gfTI4LRO6krGGoJcQIg2P1iiAqYe8R5uGSAkT/52YwPwYvJbiY56NcSSw4i41clP
raFV5AYbNkv2QUfFxnVmgS57EskCx3yLd8N+73W3SUWx0VUUGd4bugy5231T5L4l
AL93wh8BUSY/aNATA3wjPr5udZ6JtT2GcUoqU3PrKNOn9Ry1FAwJwnRudA8zMZ8B
oV7NW7l+6FCbU24BIP1lDoATTtVSK/xeruwna9/rcAlHQ63WibVxGZTGgzGhnM+c
LL1pCYdvwKD8uKc+eUCmN5po7nFSc9x5sjyiPsizyVEZ1qtK5+Zq5XIX2Idovew3
wm8ZkXby80BiLUUjuTz4SdOaBTODMtTmJLAG1UkRRuHTns39d/TS8kNJe8tdzbC3
Vm252K0f0QBq81IU6lORtl0OxMen1ERkauoz9O/EWigut4BkQPAOG0u+WJ8u5EHH
JqKWAKw80iEiZc96rDytoQXGKTGhFZJ0PgyviJVep6ZfzolheH4JH4M6BoZnFWOk
y0jrOOhaRH6yzvlgV0BHdEUOtTx/M811MivahlhfwxX0NlJFv1nJWpmK2CEv83wc
OZ+/QpE0QyAC/1xklYtykrVX2YQdWTK5Rdj8My0ia9gxkk0VZckEEUhKxVobNkOx
3lt426bTErUfQhRWjLdvRyfmuwZIeqy7pxAtFCRAUwiSTVd78PNxjbjafGBLMase
DKSuCVWhq3aWkjpt4vC6ZQ0T/wIb7tCUlaDL/1UI/NWl2M5Gm2s+1GPH60TNzARK
0mjFa/4dv2b+nOoN5jp/VUt2xmoTei5s+bP2pjGMEwGAe0BF8hfeEXhQd4npNdpX
MI9YZnbkPZg0JQVVUZ8zjWc4ur3ugAvVTOILuf2uHJRDaCP3t4hHLeMlqmDEput7
oq2UgC5CnlOlzJ1MV4gv1RN8YjCYQKpwP9SS1ho7MuuLnjS3myAwOj4p9ZH+/0Lb
WDU3uK6nEruO0ytkyuxLws58bDM7E6LwtRUm8H4qlpFH0wDXcVnLAkQTlZf5m05k
hFMJK9UVF8V2qjNO1tQ+ysbt7HR3kZq7wROKHg/FQxlybztww6Bf0TjQciKl5iDN
GAAmEdqA0Eb/dWjcZA6K2I18F+EPVWmQU/gtO6FS8s7KR3kJb5W+pRYq7h1+YYX8
8ifo5OQB8j3M8ByvcXrwnIR4/9JN+/Nv9uXR1DoCLuKGusLRulIcmBoToJ3KlF8Y
58kq+k4BpflD2L3Sam1PBF6LPxyry5ictuYkYXLfw8jB5Cbcmcw+oxICauMr3J0p
8L26W0d5XBOCt04HCMXEsPRda40h6iJZ2nzvZ8IsjnAHeOs1na9SfSXuUrCgGibw
ObG4XB3qvpI3zUW9g5EI/uz+uMld0UAoSNdBf+M7k/Lex1onmiTbSso27Wo4IOy3
frtuAs1VS9g8aHTfw5NcHjpssbtwwDU+ZycGTtHSxwSyqCLNcu09vDbNfWXHdBhr
7XXsAYc3xoUdqrWr7AQ92JvL2KuEUMYwSa+VLbRsuGXd1daMVdEffIqdzEN/SRkP
2N9AXOZyrDOUF3DE1cAyGHaeKUds0bcCqavwaUmhYIwbD2uBLZ8dqsPl8ANyrehF
gXfVAZ8RATHtJkPmwCPNJxZhoHq8m2l5kNSUXyO43QtdbGhmNJDRYar5LPwEVFRx
QBo3xNrwPx3Z+nkfBQ74TNVgtgyTIcvkFTRKYknrjolqn8abwaa4T220L2CuHfXs
fROD2FlBwxhGGWeYLu7AnBmSwI2QmQjB2h7YBFa3CFGUKKSSVB/Hg+vyJ+mChXnA
eWlTavaahUWwSa0kolsZYATc1OwjFCnCpIL+tmfkAjSc37+7CHhBYhP7iYEH9x3o
YDfRR7rxHApH/S3tl20q6TEJCfvqTfVliZ+IzqppTnRBS+gwN91A+9iASFlLgG9G
N/6LEHEaRKv/6REsFkW0aBo2QhL3BZ1kgwwaSPdmtOo+rcnOoA4oVmBHXP4bUGU8
kwyC2DPhO1jXcexF1ip+X0a77bJMB3Cjvje9fYAGTuH3WGq/pf06VvOqhbh4eZbx
lKeeh4Y0FH+vahwyucEZAuRz89cnikhXOSu6HUUNoYe2pP6dw0ZscaFacyORyN9E
cVDO1aPfP0irx43XbCrN6+FmJdaV5bDpn43DZnH5tCx3vNA4I9cxcU6XlGfj5I4P
3wF0vjZsPjCDIN/mltkJxQ++wBIH584ha8SnJLVVB/zIRo3+uPOENe38G3H5X8YJ
HO4+pU1M4s51I/Xgc2xTaUifbk+hs65580akZIaKTVhbJbuLNqrHZGJi98HNqwrc
SRoQ8CSd6Uyex9kr4hEYZ0sdpPV83HKzu9XtmT4yiOr7eoeXOKoU1Hc9bHoUxp6X
eCyJ7xNK22MsvlYVnq3hTyyN1XXL9z/YfhHZ6K9dy9088nPNW99MnTb5Ojx1/mxQ
fxLknOCg/z6bD9PjYhEDWzeN6VHsMBOhOp+wtXG+xw1ivl2eDdlwM7v9WqV6d0vR
C/agIno7Vxl+5NaxwySZ6xw/FdFJU1f6D+CMKIVKLZCW/7TuqcaGLE0IP0hhlqbi
FHYMWD22KyB5vyYG44j2eOvISCHdZkEMcYIP18RuQPWwd78EZvhadVkSVt2PTFw3
+njR+sj3+u2A5Z6XzXdgPg+uTaq/VbmIgkAoTZ1UMmgVRN37E2CGsYluDQyQ++Wd
TEUIsknQhqq8ZJLH9LWmzv32I3/wZdmTs9zg7pUNldedBB+1V4GmiQOw51xH1lrG
sKZ2+24iqwTghgMZoYIdPGvS0BbMJ95qXhIjkAr8i37H5zGmE1iSbMOt58NdxCL4
K3GFmO59oD78nxsYADvzEDueMQoSMt4OcY0G0lRz7+Lka/rSW828ik1wfol9FHB3
X1fhEl+WIfLV6K0KUtX8hCuU0PeKy2okdxskfO3WaQw05yIrD63UYt/5gJk7RJqy
lAb+3ZH9KmToxdI2DHOpXiKd9gqbLfQIHcA7UWvK6mQofNW5U95ubEoFlqONE/Lb
G41zmtqMD66DOX0fmjxWw90QGTQjdp9JFtRuIOHNcGZwrn0DbZWwqSoqFuBD7CQP
woW13M2CwusRP0RRIWV9wu1u+n4VT6zbXUav1UARglcmkdCnM8vWRIXdsixETxiN
bAP1ulsszyivuJ+qA6gWY8VMYzMIrv7cDRfi4o+FYgI7lNBGC15ipY/CQyChnA+U
lA0oxCy6dXOpoxl/pv7XMj8c9mfG4iovvpDx2//nmei3tRNHo1IJT5u7MkN4CSo2
ZJzofbcPsMlC/wjQgYkOYG+XQKRyV9u+Nxxo8IagXcHUDIT3Q0XsnYx9wjU2n/bw
n1A+0IbUVH1LkXpOiZWT67qJlp8Va8J+anNs4luFgNRKpcb69++E7HtignXyZS+k
B4h28QGWHKWJhvp3XZl5hV9jax2RE/q2YcJ7/0+3W+ENBCEXnXDuNtXQQOjaSybT
pjNopBKM9cpDs9NfQ/4PV+XPVa8jXeHyJ/NadHu1pvmSdv82Bs8Rxxk6JA1CEAei
vB1vXYdnq3BXbOsurqrGKtAATz3mkjtr24LOWqNe5ZEERMhDJjiiKErdd456mEbN
t6hv3pPETOMvKf3P2m8K4KcaVfHZ0vj0yxfgHXS+/Fwbxlu6GG8C5Ms0nzjxc34g
vqfZqpgVm5j1eMaAEcCJ2jCiBAIKAhct4E0daqJXw+AlI7C88oERSfdhxtKNAVMl
m7otcJ9CkkMuZGwMMA8u0d0yv3NsQMRT5LFNdrZo7EiaD13+EjXF5n98Fr0UXQYo
hVwSBoMG79NGHBIWSlE2DiSHJMUsSVKpBIUSwa60yLZo4fyIw/HqNr5CnJyXGJAM
uO+0GVL2jZg2YvjC8jNf2psOxbaA8B6Z0jobi2O46oewwYDO5/ZF6eZgfYuSrIZQ
/teAZKqd+m+oUOpTylJgfMsCO2VRWUgU/qop58QWmlX0MH8p1zt9Xlkij3qCndEE
zGN4uq0heHDx8LbZ4tkTNQGrPL6+mPm0ofmhAy5kR43LV0sxr0EYWBIs/75PVmFG
m8pQoMt7sYnmdZH5l28VrKlVsTBbQIgCsEeSUk3chZwE3BbUtE9Femy+B5cmIX5a
ezJ8wJbuKPV+F7pzubX1sWv4blPVoEDhXWHw8PiVwKqWd68qgfYku4RCzKq1JXVE
zBCEQAS5swjhs/vV1jYoUufs2R0o1qXzr2omLt89iezHeKyGhuuibN6YQtjRYSev
WJCBy5hHRNfAIbw+ZSsah+XOWrro+qnq6wb+FYfAAV7nS0GVNk11R10K77O2m6IO
tDS9irUxlQAi0aTd1JaxEBTXOI4P5zBjhHoI0jXVYX4/i/fECBbOXZM8ibYsOVNl
/M4R2iahloN3iM6V2Ow6U15t+KUv815HBHlj/Jp0D0ni7dAdpnZJ4ZXeluI9L5DS
o84Dl4uRx7niI3f3nPMfqeki40xxYwcZQUQVuV6qGmP4ow5qNChUe02obb7rDw2v
xwVdKcmPeVI715NK+ZM8onESyp28tjXf72+/9lYupsv9RnvrkGoFHJANYU3Y2SCl
VoGlL7q1a1jb2uvDIvZiYdXR1sOHvsPmULxwpKHcObiLLct4WsZoxUm6lA/0A0Wd
mX0d1ao4T6ypR523pPvxET0DUXI1/rgM3zTfV4aiP2E7olTf0DDccDbXTVv1cSiY
bk+UuAnAjs4sxdv6j9P05C/yYy1itpmnWotWyJzUpE/eCSax0xTCeL0SLJwwcuHZ
abxQPBSUX2mgQWaz2Eoanr1dKwB6YrAsGEhlh75QCDS9vdGsvrQXjlmOZsuo3C/2
O0x00vwBXrn669D4+1t+hhuBJ6Jv4LnClvTUtLiqqfFZzQsyk/g87iGgCTZvMiWv
/nmH3/qZFYuOF130/j6DvL4slryZfcvGHttpwnZ9JJLW+PrHXX8P78LwTk7iM4Qw
3E+uHmyUT8TQAwaxZW99BoIFmi1kdJMCg7g5dlfpCRn/0Sxzbr/HUy49Qsuz8CRC
P/E6C9qndU6P1D1NwaESJ/5Vb91masHR6L9qJAxXQmn4edrIenJuXaNKMnJydcyV
ra6Ix1e4R34dxTLwc7j/RtnC8HMyR0LM4Mp3yhzyCICM+JIcn8WgKUUtgtKvkgXg
HokX9Ex8SZgt1XXOhsjlOCj4AvASznzQi5fGNDssQFbFK0ud40DhJLAldsawr7RS
8Ycq2YTHuxIiINQ2CQ80VwVTvcl4i2fQsH0BocuejZOEyYzAKw7naRHcIYscupgN
NYl7+oMAjzkBtVNjar26z1sy+0hW6YPcpWTaS9+GNJuT0QPNlYK9AQdmEV8nXxfr
muBUaWLEzMc0jILmW068eIm1xao6VPWn3BxIdeHd3+V4q+OFo9rcBg6VtT01pbEH
xacjCKKR8Z1ZNvy25p3nIZbHKNRDnAC+TulFy4VGLo9RcKPkO/M0MZMjjxwNJplO
paxPLvZaL4NXoF2FnPyU3OoJ3WPuLlr6zJOH7f7u+ilrkXa9NqsxKaak42HO3Qx4
TNN7rt+kK6j34+Jj3N2HW4V6uAvHOHPfjd9D+w5uRdsBohYib5RPUmw9zD/ZEJ/2
Pci4AO9pfVsesNzOxW7pcbM/6LIvrXjQ/228Sj4VKZGvBYm44z0qOMXm+GHhGNoo
2ZGQPwDHEazEt9A8qXNFzaLGnngWAJA4vHITJSCI+Gqqx1kNYU/sI/JB9biwKOoJ
/A0TbZkM/RxxWBOL79kJotOau/U9OIUZuF+opomXnUC+bAtT71y57gjGfbuVSmOr
ha5AJs+Nx+Cr2yw1ijbXblb7uxp+NPLJRyJHE1ZIlxb+uc0XfJZ3XLZOdP8D0OW0
HdfjttaoLtzI6j8e8bt6tgOVeIeXr9qnIsNQ2ZcZp5RdrcjW+CQjCILMxv9LLVaL
nGl/TyuLrTRbDIGQ4O7t2w8oO/V0zpMBEludiWclnHnUJ4UYB4EArcWn3qqPjDjH
nGqY2YrTWU7gHCLOEzaXpek9c3sV2oKF9ABBTjgYmqR0hTm3dU8sNXnWRzK6YkKM
LhyeLptBHLWNvM7X0qrNhKt826O9pvzZ7oSmqI/Sl1YWZjd7DD+O2lboWdF5Vrc7
pYT6K1vqJfSIiE/rWTrev4q5OlzIPCusLM2WWt5uHr/04g/MSOkAqqmG33oWEfOX
eZ36vSP4sg7/MZnbEXUsvpyxS/DcCv7t+BLmTyw/A162n5COfsmcUCoUIvy+o1G8
H/IJX3CsTdK7I/Kdxqa/sWQRgJkEdxQTIf2+lkwdg1M6B0bzx1wTvnamI5e8rzrs
8enYLjfvYPgaa6YCNh1RvIi5oGmRpDNpaZK7l/u9GI5ZIfRV8UYqeYIoICnTqge7
/iyh5U6dnm4NIxgFvGsJKyYsbDk8ouvbM60bFNol6hSiKPMrZ6H/Eh8mn5i6IJoS
pZnEvESu0zG+ZsBzLJjJWtKJcQYMzHPjeGT4SZVS4evvh+GUT5ktfVwl8q4Ob0uf
foQnXpvfAPyZN3daayLa3jNkj32Fnhli23BmZOXiqLxkOoVxEelcipqAnwah3Piq
UdYUZj9rGXTYSVzUCKavKG0/c1y4ywv0IyMwcbxkHrRxkDVYBlk8NAEfcIjDW1Dc
HFr+mqV4VZc5t/7dAexXTU1DY+oyJhE/GrPvtXA7o1iK3ay0P5jnHwi2fNgtBGrA
STQLKK8JrKcjMjtiwW4NqjKPF2VwhwdGBdVExzNYpFUxU0CspScBXR6zelKF1CPr
/eLd1ZeTO1ue4MLfoyzTvSsITCXPlyYabjFtD2XP+iQow+wZzQYxBVL1xpqJ/XY2
PRQXte0qG3lW6Uxl6akxqQGRXdrDZCjJNQN+ggzcmVYeV1DWwzhQiu+/IvM7hNZ7
Ws44vRQDxW1yXOVxpGxnHraz2+pRq8bnqMFN5Vs0E1V0CzUE2PhThCjDpaXKTh80
SZ3Edp+x0Qd6ggC+h/WYV4gBItPVlzii5wrZucEtc1y9QqsTSM1jupjM0POImnVe
WFlTecdVBhsv3nuVFEr91K5CHJ7oc98mBFd7Sh4kmIFkJs79SDwrXhWqgoEv5My3
2eZ/xFsbzdlBwpvXvnBmeFeCxOOjJLCl38+AbdEpNiZmRM2UqsbL43FXk5q+IaY7
1Y/M8pkF+sY5eySNGKTnRvivimJkOZ85R2dxNSMAW6SQriP5TiMe0ZP8WieXIcIh
jkVIKoWSflKcscVrlhifhWHyVB0+remwQBW50kbC3VUD9fInIaEwtAWdiFwADWQJ
gOXGGkmbKTusrZdvcgKhka1KBTzTWYM/wqqwZZLNcWwLJvJUxAAmTN3nS1LNBIAb
qYo732T7l1IErq1ehBT1PeCSiYYuc3DLkcCQNp7DL0pCbMbZ0SkwN0u7VWXikyHr
LHIvwtmyGOtA77ShjXITDN376A7RJPDtj0qCKHFDW6EMdagL5bG6v+iol6O3dJ61
cuPQnf96f4q7Ad88GvzNjQeVw2GBRCEeA1rQNuqMXBmaQxJx+qLngiVAhppcRvGi
bbSMDG6ik6ftDGnkkbGucVON9Yz4q0k9mHPo445/H9eVALGJIhjnAaUq/Tfll6dv
Frv3EUTiS8XwfvmdMqwMZwBhZlgVPWf+B/lxqyxJfpxTg7+nBMfLqfa1CRBf0km0
rXIc/QVx79LfZbUPU9bMfz0KAsv/R68+/VIVH/ZMTpygkkRoNH0DgL1cwlng53jg
Qxq3DxS4GOY2hN2XGxlKYN/wpW8XxPeSYZ4PLOnFPWy1i8YnGIomIcBs5hsAy4MP
BKUmiY2VOImMEhmXoferD1Pm2bo1wOVDkrbVJoS2E0uw0MaeUug8n2c1usIwHKfq
x/sm90rAQxwmRDuFBqUis1SFHuX0CY2f+N3ExBcAhT/CoikjMAxvkbnaOaX+nfS/
sM9Nzc5eZM0N7B+TDsfKGoAV+VBQwUU0wJ+45iD2yv1locPYlP/eQF6o4D5LAq1L
g6j7jDshgAkBPQKTsfILWJ7gppX1zoNGYtNBF0LS+3o2OsB9LqWsZBuR1fQ1qswe
ozd+fbTldk4xx56v1pW+xScZNRWoK9cu5a7Ozjyp/HYGg6naeYpdQJTCMPJbCZmu
mbKj3FISkVzEgF1Px5OMyOyxb9Wh5cRs+IWVMn8Ub0yaO9atT+XCOd6guGzSJOWh
zzws395LLnoYwmrZKWcW8J9uYWfRpzbhAK1vjB/LKPvWTwFnbMEhBzosFaoDn95f
0a0XQGtmDVrHGxxK4niBqHdDTNplhzmzwtxyTzF0osxGGgFRwOhYrPPQX8HnfcZG
36GS2HwUaUUg1JFJWlUZ9wH0AGXrhUqhUs+A94p2vFr/6zZeDvljyyHNqFwaPavX
aMO/G6fBv2du9o1mBhg6RO31WyN+Cp9ZyCM3U/xOVbhYyjensI0vJJC/7l8XwJWJ
y5gwusQw9+71ZL/y6jRtVTIAuHCcpXpfSc4HGbq+7ivByPyBCLMCxHWv1Dls5sq3
RUEUQGEXb3XlViBQ2LUBkfK3OO84MeFnq7+tBtkxWFh7Mrk/ODIPpRnTworMQE7w
YdnzwmZePoOYl/CLsYJVFE4fMeNqX8BSjXDlgLzHgjgP2i9bWwHLzZv1M/My6gvd
scrU8uDLNBISJzScam7oxgZdGLhJ6HzAH2puZ4Y8CZhs8o5uVykxnAaz6x2xoLsH
d9glrCwZdNS/8gfUGsmGcdPyfE1dMczK6F1LGNlcuinE8tXtcH+yEA+ztxOsX6ie
ulMJh9Wez0i4TjOc7+hTgcg3fcJ+WwUcdz0Dodj2pHYdGgk8Fd+HXuwQQGF/MJTV
t2K4rQI+NzwklvPkojS+PAukHCrcJgUbqWFV1ZA0HKG+8vzdfBTg62yDNC013r5d
PfxFF++OQ3ja3xHfVFB5YvrevZvdP2FRoGjG8/xMKgx9PxGGbLWRKqqh5P8Ge7fn
kikhOlhe7f6Rcz1+qujRD+cnd3bSXxdCISmHiNfZStvQQfVZ/eonP+eTkuSmMqlk
MSP124RrjO7PFpcWiZrPdTZleXjFq3q5b77VMi1iap4O2cv45YjFGnAHt09SIX6g
F7YskKbpPr412GQa8m4ofwABLDTXF55I8adQX73NVVLgM3qF0nTdcslVEJMRE6vv
SbeeEo66B1PrrsWugLcWcwKxkRmzeiqMK/hQRv5p7H7aBwVIgYoivGGEdqEQ7EEe
kZQQlWSZg+EW2TUGcm8SqSAzayj5uklUmAx1ujN/LLuTesMcvWjR0F9DEjVglo7t
GoHU+f3MbNmOoqIaYWhFXjdjkWcKf1WcYS+gVtcp1pgL9DkrRPkA8d4oh6eroX1Z
8CvKr2yf6U+2oGA01dWkrBf5wb7eEAY03da2Q5dNmpwrOUmcDGqCySFFRNxcTmv+
+cE+UpHvcyvN0BSOIej4CIhzOLTOF+4sk7kJt3EFOFKRwBCUuy5hgklcpoLaC9Tr
Ky19bB7sKCyoVhRLxJM/m4NqTEFTnIER1eVm5VMy8Av0rHBzAeB/MJSRpx+1g1Of
yedCFm5WWctZL6Ntu365r4YgDGaliSTJyGoqwAATDn13NQBizE27qBbswp8rPfE9
nDmKUwSt22ISjPoAoFgoOzlrLIwwULqS+uR2VCyj93gNKXHG25waOZ4j0A+LvcmL
W9wgpj1p8KC9Vmc+W6cZwz3RlFasBaxgSSSiqXVAUyOYM3BZ86RyVUKGYDp9KjHp
J+gNQv7V0XOuM2uGVujFoEZtMvuNBOBWFQ/tJbQWXBAXo4aabiIMDykA6BqqScUS
Pbkvk5q+ASBdzy4d4vbXyNzU4qzvuuIT85pD+Qnq6Ituqw6buUUPOyrWQUh9D6x9
ycC+oZnI3wfByKkp1dzuNX+Z8rGNQ6Wq8Ce77u4CavZgJm2ClXkAfB+oz7kjqYPQ
DYtvtobyw2VESJqqRvP66KDfoUH4vCNzMIv+QS/FstXbhVYhAShcJwlnxC+/nwEv
h5b/OocvBkSIcGDkhKPaMo3kosrn63TOVOmNKBSa9uXf7UF2Nw+uv/dcj8AN0yF4
HxXDVviKYbJUl5WqLA1ysrtxa0AbYnIMIRJfk8zuiJpyMXdKB5p2rvr/0kfeVNMx
G5xGheaXq5DP7PolUTDkP85Nw8EfdZJrzL/Yq3Jcrj5XllvFZ4TTBae7UOUzUXQ8
+WD1EGxOIRCYMhOiuLZDmVLE8fT/1vCsTEDHd+UG1rZ8bbyfSLAirB2Hd5PDGVBk
8jU1ikQzi/khSvkuXD4Zz5iwHhhnYRSJ2M5KrsqRmsSGX02Qnk66bNN10yUrpmQK
KsFnpSLA7rVp98g3OTvXWSwpmsEShdWyK/LQHGETrxmAZee09TK+i++z70z8bEqX
BDWA1MsjX0SfASeVWp0n9/kdM7YccwQ2HXt6IzcpFxOgW82j2194QjGYEBRJvOu2
nPesBVcEzsJ11605xEYc9YRQi7jq1YNLZC+zAtoehal9Hkd12oROwQpS62HmRQDL
FAXHL0pAXrvNPUFmN4uG6hlxwYIl82ppOXw5/K9/wszSgHGOjzNODiKNRhB4xMB+
bUdCGa+vC0SsnXV4ms+hvPTpQHgd8F9jthSoUdB3cc0Z3E8+iHqVOZW104B3rGtt
VUNmfKfLblPIuhTc45hSSp5u9/1zv9Qf5ajH1Hwb6JjDkU+TswZu3mNq54Q0do0j
yixOWBqbb8aqO6RE/N2MASXmiwjdgglznc3zuMuYTs+rorB0o1kkSkGA+3HDtntu
SZ5N0fsmfrIOEYQbXCCeA1yB9fy10EHXWBq7al6HohUzVEY4P39rrJpBvPzgasc4
Ud6Q5RA68sooYvYE/3uyXsciR6DSKadEQpC5u1TbTXWvu9Ye4V3Ipg6WCdlrj9ly
pGkxDdmqLaZAoUjGWPvO5j440nHyibWCa/coIggdsVHC5qBhUG3xgL2/XdnwJD+Z
c1t4RF6t1Y/LmWxWJy8nekk7oKZjWsXPDio/l6ENcmz9wYBJHWBk6WV8/ubVHmCP
eLJwFYRjZzsyn5jlE9lyMcOI7sGfdha0R4x486+POKZPABVNPVpCMq9UhHvnpaH2
Tm6HEt4iKUpap05Utrii8wB2Y7wMZPVjTa2oHHYs34mj5ectLzB4VapSQGefeLF8
cjk5UcG8DTUYPILFJU5YFGZenncgVFJabUP+e+9tDZdAdVX0Z/td8FLmsss5vn7m
OmIjKkuSfe9gX3GtG7K6jXY9y27FwDPLV0nUkBPvK9mFtLyAP6AFu+snTkARtj91
cSszxEqMJtRVUGVOJBjN4R8wnphZRkz7QxA0zX+u35lydQ7picnsp+K6uXN88b++
AabBKQwkdWAl05M9HhuuLig9aclQzJinTqLg0AgENI4+/zi0HSvAaS79r75d2Nqb
PS1ymecihGsqYgHKqmKDiSfCIqh4001JSkdjexXjeTc9qydIX4z8yjT3UUYgl33O
5KSg+MZ3O43x693jhZOK3xuscU/1u2lTxtnQuySczNlT48C+YR+T3TfrR0ihplgf
7Z3E13qN/WU/Io5tlxgmzJ4M2ddeh0x1+Ac2dVzd2w5bMsvmsioBocMxOOtp6wGt
gR4/LGfshOP2PmLkxTdmd+7Idc6IVmzpdaEwSYy9O3igF0XzAy1AxVpDq/jSi2ol
9s+8177C82n7QqU2jB3U0OZYscAqdNDMicHkHmM4rtIAGRsukI1QDhAlRvfdte9N
9nLrQtRRX/HBSVfQFlXYs7d7x3gX6DMbQE2Hg5lxjLvy+F3ZZ/UrWo0tMP3q5dAq
JobVoENDd4IHd7ndIA8xw6bzMGgbF5FVDNznXc7FDj7CHXoHQwRjAGLWBlDMDWYq
he7v012CvmazDd5l9qrLDt4AzNWcHnoVKyy1rQO8jHtCQ2U7QusEHs7BJiWB6car
auxLznMtlry/uuBuIdC86CTfj60SmJXMPqcQ19mMiORuxke0cR/hRxS7p32BRP0e
kyo1doJ5q9y3ozD4cK4OmuSwSox3ilLUTvqBtlKR/Mj60Ss23WOrUPNRcqPI/mwm
Ahnw/+ZW6BmHsXwhXZdnmnsPm+dJ3eiFPjpx5Vf2Heu7wMZyWzCwXRSh9hP8OOuD
He0xjecdBclwQxXYfN4afIrgkQS2e+BZrmqsZBag896X8Hq4hKqkU3JUkz0W9tIA
OALASHZAJvi+DLLrXvAY+g/0sClv+A+Z3pdO2WR8Qtxds9zaHhlzCeOQgKOpkGaz
R9EMi9ORtB4PYQFQF3neV2NX1YPQMEi2Zdx79GeZC4UPxYmW6/U4nctNmFBeJE2Q
dTrcRVAzrFRRiXulLTSsDE0e4NxrFo/46uRos4B07y4llea2VBbW53zfrTr8xI6a
SUWen7xCLSyprQ8RGlwnk0PfD4+bzz2ejAZm9BDeRb816e3nfHK2PD1WufXC5/jD
1Iu/QY+rCiVyWzLCsEb3Qcs1RG2g7hmo6XEjbXim9ZSPtzbpYQD+uNpw1svG0U/h
CgFHHreg8yif9C2keOU4ijaxxfkv0S8pKWfdYdg72ottoaEL2XiQiJsfR4LHVvi7
X7MR5ZrSZmfKkwi5tvQgHOOVxpzNsxDuKJ7bRN8ryUPwLc7z5bWkmHbRlgPlW95C
kNlho8915KjzGES/uTx+vyfqagHFQ+CB+AgkPsfY0/SFiox2sB1K49zVYWBVXFLc
ny6x3kd5wRnCAgsWtscRYq4Zuc2YiQE2A3K3wZYXYV7OL1lrbARZWJtQsfbkAcQu
0huXca2PSvkVvsVt2sZ15xmAqebfsueUbVxFvPKfoFI9JlSWN9Ncb56JvsYoLfEY
OTzEcRRr957XXv03mgKHSDpGXlC8sSBRkBVg2d4SOrVNirvczC5+N4qkLzsk/MsX
dFFzhB4I8b2/dpbrh+a+aKiAph8N3CN1lCEAFLOZn2UOc1gSaEwfqggXL05IcqNN
6b+VhhqtgjKIcWUOdCtjamQ4fvz+tueXtFC3TSm6eVNVRUii6teDNQft8gNPdKEi
8alMN74jGnnX5XFKp2XPmlqqmh9C8vT5SRHKz2Po4OXfXNrHI8NCCwXIIqUsFaAJ
vpBNKK//fLVHYooRn3BN1vjTD5uBljXeABjRBYIRvpyrgNtGWqG3Kxkdh1IEt4dA
AjFQCP7gmEFOMndT9MdK7zd/eqeIIMo5/wXl3F1lNcvWCFUDHlr1EopQXW9FmIih
25Nl3Y3wUUSRHlzZ8OjDVJcPyo0CnxM+XS6JCBjEgEGH4WOtUzUGieg8Dh4fqx1+
ZD+nb1JwBisdO2X1IRqavEQ2kBmbLl+wzQeDhrEzwhom8UmravMmI2JzHeHYmNCS
c6Hc5wFM+r1JWIrFglQRKfRu7+UVbqf9boAs8JZaNtaXPaZJh/pE5XWJkVBLT7Iy
ZtGUerZQCNGWxWRM09kHAxOlhNVFrotR+k9j0uNxFaNBRr95wOaKO5HyrY1AHiRK
1wSo1cwGjdPydnW2JIOwxzLtSFYLzcDClRgpzYL9bAoAkok6YSIe0eSy2u27RHa8
3dfxB8+sVm/2/Ed7i9JvaUZoo9EhOSpUfV+pO1JQVqq3FGa72jBoSX15ogdxsDjY
3TCrFLX5tMuhrkUyoxnHPKSZNeQ7dtzM9wOXr9PPU5M+4uM2dqG36138Hs+AUfhY
8CzQpu6UsKMj31sdx0nvU2Xkz9zI0uEIuEPDSVnTXdQU/eOk2Wnv4p39GJ3YccVt
vDB2FNgHe7at6eS/HY98IMcL4S0pJt3VPibzTy9Dol92E0UAYHgIMroKdb/PgyLP
vYiXHLA8q9Gji2EfSmhLJmaKRq0zQOMDXP6sxSjnNx7tV7qA0qn16C4gTzyTJ8NP
2+tZ80tx6uOM59dzrK9ah5RwPPrCfxqYtnOVhHx+AXXWB49yE0AXVYa9aobSjja7
6CZRhL3XWLQPW6BryrPfqArUdKgcOpx4xfdle58cVldqtUssOYfZgzqkjnNYjpRD
SDHjHr9EIKwUIVZR0iExage+gZf70J8MkZuGWIb2STcNBdSoQbRckMpD7xDVzvaV
bP5bG3wjEB/soLwGYvGDiOSylUBPpgSvF93zGWUzRalUAZF2Y6g1ufUkyB78xd/H
Weij4uHu/lWPL9uqm/CBS24EcRH56iSuYnBzu2TWWJBsut+ve2eY0htlOZj25XAs
0ip2r1N/zyfEIaBRsKnrwbwgXxawuNjs0i0wj0ML+yS8Dx4snOmx0iqd6tg1SAMw
MDa8ZBoIbiUGZaDyJmiLviRuUZ0gWdN4lm67qFwnc2Msv5FBaFoJJpGYEzSUO0rv
+uNnUmj07mBIUTY+J0hE5h6aqi6pSTIdOP5lhwHuW5fXB7FTfID6oQJDOwAcxmCw
6aqpDKFhQcWhjk8T7WXxwcVKp0jvKqmj9wACYCQsvx3uEEHmor0qFkdkc/b90fUa
8r5JYI/waZOl5tuUCnTAznZsi2CAwO8+aRghnrPSoUJcGR+kt1pW1D3Mp2wXzOp3
GQNKtBCvlKeXl5DciDsoOYLBKxEwJR1aJQ5Atg7qNdlnURQJ5gs/XYCB3Un1xqzy
X3K0uepO/tZ9yRD9F3im2hiX/nOD3O/UVKspHwKhoV/+YUGYkPDqwLmHTveUY6x2
Ivlig5RMcNLXkviCA+2EWttCjHZd7uaKhvqokX5dv51ilbpjWG9Wkk98px3YclMv
+/NwymOT4JicMGBwaqqqtZUPnFbwAN4LYBEEVqfZkzClfiijj1e7WmMEAfsR8FLD
AJCtrYCSDAlAIC7LwvSnw6Mdmd2bS8n+Z4OhZjkuHGKggRErOrXhDPaUCR/agHW5
5HWLlxv8xptezcOpuJoAc9ngAHGmFTbUDoxlV5X5oBLnhzBZIadfiMsDf9GI2fRw
JcsnYcrOX7CGQMHCzgJE3XpfotXejRJN7J7FSOc4KVSRe8mvXTkvdPO8JyU4incN
PekZoSgC2pn63ZOtgFEKIK1GhiXv2hunhIuKx6ff4N7MhkIXsapyXqgwvb8z+5O0
HoB3+mOq6/H7LFYILekZOa6zDEcsBv0XfZBT/SrKsZgntLUVTFtzc03XJfikMkrE
9lCgQ+pbiQPFseZmy4NFIShREYDmfo8etZ0IMJe9cfV6XZxFOk1FfXs2QSR8E31w
LlSdS5QaOwegaaS8x2rLvPlhqdhlWg/JDQGk8nO+dV/axt8z/P60qoQhP9Gn8YjQ
CDU6jfgylXtPYFB4H6JPuMn78swJD/TK6PtoUgcPh4TlSVlUsVRrTNVbhRJUAOgy
UQDAsrGVAEv9OnF8uQqXzWPHFYRdNntMH7UH1/MdNV9+IrUuSamVUeiH83WwcqTs
FG5I4Ic7SXsVN2JEX1zS2mSGS6J+DSbeV8imwm+Jtpbm+SRhnISptzUiya2ooImg
ZMnc2rDFhW3j1bMcgrqzRpGRzKJqSjNC6xa9YTX1d043AGgPpQkioxZjM6l5k6Q6
/tKwaZ7HU34I7BtaOB1jN1JEBgqYgaO0Fwven54l5ICqaCDu5Y5p5LFDG5PKTdaw
d0YkSoPg0yNod5DuDb0W4IYiJU39HF3bU2coq2a9N41oHX5ja7TUC0KB57M56ERk
XupDRSfeaunwmQfVgmF3sxm4AeLj7I75QB514tClh1SlMYJf4fcCFoL1+2pbd0je
BeD5+M4SNbpRbtJRqkp/ubboBY9rkS9x4Xf+YhCNauEAiLPj+Vt/dkOmY+KGWiNq
3Q5EXGnVSHc9Jc2uAV5b54a8YtVteOP+RtNEDixLn02qjZ6CKiSLCPGg862RDBuw
eKl4hBzdqoOli5FCTjx0Lyn/3Sh49oXauFX9HY5I/rHC2UrNG7T8S5i+FQW2Ihwx
P5+xzO70wPILOlhBGROam2k9pU9N1HFx8UuxQ28pXGfHPfpr2iaqdw9c/zsfwXCL
QwXw0X9rTv0kCfoFIEk0WnUPfN2KpCkPtIQMV9XByxvI8eark44q98jD/tUMtRuU
9uP+8WuHVBaoHhZFUTpNGHZVodZrZtxTjl/F1J3uwVoxzc/9qUDPqozTeNRW858u
P/wjUaYNNgLuhhgTn1ky8lc9eYuoOCqqCenGdlmVBE2i75sEX8fNENNKLx8g5wlA
4dPwHLuGyYKi91qaf7ZuY77debcwl789C0E3jGe+w2EhzQoONA20YhCaGoayfPqV
QIB0W1fJM4FKtaCpdXUUb0sWr8QrxnctslhBKx+qktcCbwNNCSIGH01u9D88J+MH
67HvoceHmXVY58y2BLq2Gqa4uWaL6ElGIMCjySitoNfVa76K92UIGkFyqoT06KaN
FsFku6oe5k+7qS4yi53LvZJGyyHVywSLFGb7Yh/PaxVeAqrCBd9ciZ+DBSYD+5vR
8qr9rkF4a74mI0PNcN5c83B/5r7+c3vJdQHpfQJWnBQuYWxacvG6KuFl9PQfWfPO
UqbMiS94sfadNKOlrV4b+vnpsnmSmOllXsF7IHTtL03cF3mUW0UxuWBTBXrocRR4
YXJxxA0+RDr1OWLTUgyTx1ix9NdvDDatA9/E7rkAxD0mEFRW6AOYK1+id4Of3Dbr
a6BJdsH+AuWvzQONc7ZFazEURgoxgtPYJgfGf7AzQgDdgswkZqoF/kZ3iU1Y0T//
g91wjqcsYcQ5RyirgPsyzE5fIkt3+0SI0cGNVg3WCSQ7f8RCnCBOICJESz5h5WDN
zfcN8D4on1PcnxccejiV8+o1O9nxGrnpe0Pi3xKqz2stZRnoKzWABGDLnbE5FNHS
YW/fR4I5OhuM4wIjn5IDdiAU03NvptkGebPjyeo+QI0wkds0FHtyE3f7bBhyDk2l
H88nvwgN3yBG0Nm7gek89QITYABklvuCA+acVOJUzNI7StV3z+dJE0NzGBaw5WNP
wM9jwtQ6jXzugBov6Ny7ambXIG+RKzHHKnL51sH6/fv98mp8Ma4/tjC7JpwzbmTZ
f3vgZ7KH5plkPCueOSIcTGE/HJQ5ouRSUdLGbALJiQkPy8jjn+oTRBY9U5RMZses
gaiaJ78bPFQPwG10CXRqlQBJBFhFkfGSFzvAdwcxu0TAxATFrIRjzmDijDdyKQPH
ZI9bJ16Bng8k5CiJ4Jvva4inooF9SSvhRn2xy05syK2uCLAybdEtuDDK/J5LJzsi
/xzYmN+SrzG+K1BmpwXqfI3ujQcUZWD8FYSq1F8UYoFTo2UM3gFESYBaNAKtuMWy
MTopAocWKjAcvDaOTRLAsrECgVEYBm5grKwYiITgNFAHk980RucAAQeoYRsyyBRK
K0JMkCXN7yi611euBSV88nG5EXZPRsVu+I+dd7jyH4yJaL3A1u94GUTnqIJoh5Hr
m0CvC5XvE/t1zprB0zSTKpi+Tsl0pWgec7yQbREi9CvvbTt/DwkgokxEzpRsTDFq
7XZNuZZFIZIG1Ug41m9BBXZDd2CA4gsnPeplJlfMV3m5nQNK93KPNkG1fGjGFGm5
RH9ZEMo7VaqIspP0lFlVjI6Vaw3Y4RPE0aB4JjBteUaQk96+eqYogNfuRdYiA3cE
J3xgnJ2RFuK3fYKaKvrSoKKDQTtD0/Y8nz7Awnmi6SAJwSbwfuuoVfR+VYQpIZhH
N2grIg2VXmG83c9RhI6wXGQvej598PgQYjxur8a+oMP8pbtRHHwJIQqTDUKERmsh
rBm8W8svvFsHf3I5L3XC3u+SYzpvbpS1Wpkzx0FiZzSiLAvZHA2/8Xpth6eHGTYB
zcfB6A4a2pR3u+T//hbuwoh65dQp+bBCsXXxGP5rzxKl2S/WATiafF92MF8eiGP3
cBNHSf6cABbxkUWhpl+IlTDI2NbuJH8AHpPAY8wsBhPstLIajWd+PbARyebCAiMK
3w7xCANToL8IKH9N54xKG6Ih56rJCoHst152BtS5Qlr5z4xJzl/V+Rz9AnKiAJ/N
DhX6yR6LGlfJ6kRIjWVjtOWRY1vXF+vwKJMMcZvufpwJ5tD8LWAM71ZDTnxtlVmv
f3e0GF+M1B/fdQHQxTHRaZsjC11IJ6A5g+UOhULayuUZL9eICJnZj0dCbXj1Lj8a
GY262+ogladLEIkCqa2Dwhaeq9guGUlXny5AxsIGnepDSYvgbxCCWBaTzrvHFugn
6OmN/MJEhxFA5ilSX77UvJfe5AYlNOZuSxlNiifSi56TXfNpmqBh1k+KOzIBeobd
XsOqLQswFhcwkYBZVpk5jtWwu8UDNJa4wTIIH7SrHDAMt41monBMhgt2bx1YLQsW
Ua+1YreOkjErf+kcp8xrHxHtBbxmHh/9f2jpy0MUA1D6NBCDwnllOK6wmYJMp4QK
Q4amTLudaRAGRLbUxH5lP92G4OdMUDwrgeYyLFzGHlt8E4dwKk943BoU24g5HO5j
OEqK1bttjxD2Ocx7LP4ogzEsyi0BKW5w+/AQ+8GXHXB2z0s5m4y2ako4xL4Prx7H
71Opq9P7MGL4NuwXFtqqgNFI+YiV+dOhDs2QFiFXjTCSo/1LfoghAWVQAkUuATUj
Ay0ChoKvVhZcjMwjWSjSIR3PVq5Jd/P21s4Pz7pjyQmDHKY7OknjaUUSGnN5z6mu
MiTxpZw/TWExr3I/U259CXpooeqI69LSmvOqFddcXj+Nfm2S+A3k6ehRqmsWTXPU
OtdvIafOFQXO5j8BqRqEXFOX9S4WaWugEzz6I2Q59n5IU8q7ckb1DwyCO8WFSUp/
pZ1TPwSUTybhSb8H8UwDETeVqj70ZlXFggWkAQq6gdHuE8VffPbt/Bc/FO10IkK2
WSs4EoDBBgbBCYonsR006Ofky44RJPJ7wAsBMZLi6C5Pwh3NWb4va0649aCVqjby
V6hgSeglr9egWPC5QI9l+GblUiD2TBsyKD+keRtVKuwN/5UXMXRuvIjgBeL8SS+Q
zDd/bdYUNSXskqNUt3iJBdz22hLMfspH6S0OEYNjRifFDAnC6OoXVSynLA7uzPyZ
0XoY2ht9V25w5Y4siaamHtJY/bOwtWdNYsLfLuKJP5OzRsAVzjVrEMv2Fk+GxZsk
ED6lwtMXzQBtA/Z5LEBxh1846nBZrbtrsiCEt7MKZpyRyMvHsIvoqPYb9dkgY3hW
Zm4oOMSkSPO9QnE1D/u2xVCdEjbpbrO8FZQbd6Y82Rjpa1myUzkUijorXlZe7YDI
Cu1da9KWXzpyAy7bTjC6jhYheL3xu3Aje/MbpYS0xFxxmRC6X7hRAGcvdgJZ5yk1
A0sdUVhcVHkWmfAJuly2LYpkNEv8R/yP9/aygMiyMXTrvepX+L+J9ZEz9YX61d9s
Yg9cnUiYTQMjcdRQkO3ddsH9aw2cIqd7/WJzLDY73cgtDRUSZOQFRJQiI5bisvV5
ITS7cmhsduzJ+i2xEtuRWMn1F0dxpTPuk8nieOJh0MDPDBS0vRAzIRt9vE2Bizon
ycSEAbilB33lljft6mhfcij2pdZI5BCymsWLGUC3OgSQYL+Eb4kX00T8hn6icROY
ldYQNzG7SzzRuEA0W2YBDLwTUyEypGl/5uWQQYbyfx0XzqVGTELvXr2xnMVwKVeV
JeJvsZRm94Ws+0St9jFOeeUuxFVlv9T7SfgsMbrV0GrfxMyyzz62U58+FobEYwDy
US6TbH7a4NC3JV5Kq7jD2Zfb7J3xw30091dgTcvYiqS9o/ji1uBVoPjcPXKl0A1L
pwfPGd8mf1PkiXqvIVqe76AtXxM/U7lrOxDx8HP3lzCOn8qkgWEP1atSxv1TSjZt
zjWxs2cTb/3c+Ln5Sqj6Q3ghNUzUP3FHr0TKA+jmK7ODNol6gpdM04Hr2APxUNrJ
itZttAB1eh7LFoTeDTCIbK69zVmvviH84ZOidiMizo4HeXgPPM0qaJ9BnXtw02ts
EYaiHDF4Nswfb5y+wRy8chkH0t4gGx0my3NuhMkQV55pjQwb5lyv+O4apJ0BK6VO
EhLGOJOVxL8+oTcuE+Xxlk6BniPjlTbdJ3jSfPjCeYL0hkRMvqPS6RKnS0h8YsZb
repDxzwJCxYxxHIXoBqYiycSwf3xihl8AsAHjNc/WFNwRKYVfPdt4L6tbfjmGHU6
fQqwFvE7nCHId8ugbX7ELe4GCel/IdaNeXSucOJhHomReeEnZaGpjl2M8vblOAZN
zNJr3OsnQyU06p7qw9B/qyeNzS3nhXFfxIL4OednRlsehz07tiXw3OHezyajUCiM
OCUfurPieWQN9w/EzEexuraHt64nQbAoYqTJeIIbH0CoSjlG8pFEZ/qqBTJDuOih
gaQ3vA7fuq4flR5OyhhH2+sBGBuqvcEp+oLCCCgWBUhpwh3IPBGOokkTEv3jHm6h
lIXMIbE49fPfC1gTIdV6WxN1SOv1HvhZr/Wzwr8XAkmrI+UrEu4mKNtI5fsPtpov
EBUGz83v6yHjPqjm7TuE8VFwN2dqyqKXIAfOQmRPTREu2bLvbYVteliMnU0foFmS
BR6RnRPeJJxfuRe4zDJNoR2M/s5wsbbYywVI6ugZw4CoIp8sQpomPEykNZ4buFqt
cM3PWtQ9l7ulhu/BdRb39Y1/YtVJqLLNsKS+1jbzqFGncTY5oCqUeFvkl9QzDYB/
SyDP4YtULJ7gq03JmU7KQJ5BsVfSCNliqhY0M63C+FApD9r7Eb2PjX8R1rdFu5CV
T9m1YiCeLw/0NOrhnaCkbkyMUPCide5BoffcW/1GtAbOEachV3FvdqH1DOxmpR2u
Y+dES1SUtcpyIk5p5+lwVUsrd4TMLx3flm//LzP8dA35CUW+g4/YYKwQFc9fcszB
FXn5t2ifO2RiinH+G6UpkxMR2NnIzYiWS+ybEGbskKA5jML3Bx1vKg7tNwvl98Mb
QYfeEBSk1f5MsUvyLF2t19yrqR7Xn9Y+/jSJpL2T8NFw7YH5qBb3nnANsDRk7hYd
uWYcYLnnnEvevxrdAlqXgk2wByljJb/q4KY56k+ceCfVBC3jwbCFty5OkjcX+1Ab
K6bLFlWsYY5J23nvz+SU/r0zVyPoaMg3oZHLDW43I2LUDLxO036lOk5RJkGjMV/O
c1GwKPp2QMN5TuvtqExaNVZJbapaYLZbcgIDfZIxKh9X8HC4Y33BJlBmUAs/9PZ4
kDeitbj8xprJ7G6WPDQXuja5i6ouNiNQFs67OlJ9Bo6bKqUXETAvWJzEEk/d5W7Y
U4GQy1O97HmSYCpNgLpOD+i6atyFopj6rJujrGgTicgkegsz+hHUo3/RVC5eUTXF
eNr4J7WT9eER7AD82zV3QmxJ3sXQV9kTNXlnIk6iu122ss3TwUC2WqvdnYw9IAhn
GQGVltrE1ylnsCi2GRReaEMkd3AapAPSlMetdM5cLtLfyU0VcyVkslImmJk19LAd
88TxON56BTLaocnj8ldfLPqzka1yCnTeusgk18+A33Ywb+mIhsCvNoKj+ym5WlAy
gisK3B3RXW5CLDy7k29rQ8mJ0y4r2apEzwPSkFFXco2LLhUD03erWii7vCnTXE8w
9mGk2OtS2frJgJ7Yhdy83/nWODmVj9VwRpzsFdUBPoBRW9V69vEpOj7H0Iy+B6ze
LsxfZNDkACg1dshQ2bm7t2nx9xVkf7+Zz1QNidmz8N3txxyrHJaQbVadOPcm/U+O
H0vTu5LhLNsV2IXkS6g+6ujsAP42mGkDJ9YSlDnnRUR386U9bhn4vIoUbtmugjtc
msi1wLlopyCHw9V6fLQlXxHX3okoS4nlkfdHIzS2ZjIC2dRdKCGuS8LdHVLu0QuU
GnoD6PUG40h17h0IgI2WL3l/Rn1wesRlT++Nd7zdjZTlSIjGNRWutmcH8JRBO8kg
0W9gkd+gwnsuIt6NvqpDp3rCcVEbaU5ew/eUySx1UaQh+iFfwdPCtLbfXLyapJmN
IraAQSpYSIzEx9M55t/cgNsiyo+/9KVf2AdUz2ISi4fVvhSOdoKDWqw/+icdTFMp
mlQdMNs55IWUoi1tU7wp2p9xBqLrSJcAIhJfyMioDN4ZgOf6HanTgIEP9ECy0yqG
QG7TJRRhvnjCQ7L1NiLptz0/ixMbMvCw+K8oVRVeOFD2uM4thrS946M25h6RQqAl
2aiv9c5jUWjjKNm19ZdC9UUMZbT+b82vp/f9iHgQrYk+hJFAkuVni0RyYAqH5A/y
3mkmx510gQA8+8sW87S9YZzQ5SKTWQIg6NIkXZ0pTbMnM4ivQwLNCkPanlYh4rsu
gwmhBG5KCeyI2bl+1358hmx5naT6KPJQ8jbuFhlPYSqxVxeJ7VqhzlxbRgEsEc8u
+aNKZ1rqmiSuu9IBXVMlnvXWzDfsmSdt6UcdcrMb32QzObCymXDRXAiK2eZlgFxJ
TU9ARzenWdRebZBUaZQbFKjnjhHrwIqx7+MIVhOQpd7MJjuHQhAohe/SSpSWUZD5
n7e7WEtDQshJ+z9sQ/v6WyOwE+XXo50u58/FVbKaSVHBkrR486p60G/9hxvK0nwM
fHpCRZf5QJX5WxjmVBLEKoEPRqAokZQiA1WBhjXYGgzAG0xpNlsb3p9xVnRwZquQ
KP2oQNhpTjVoCN6KvoGeFNoAhuXBYqCoIj4qFEjraFS0E84PSzbnWmvaUqE2LX7s
CP4N3EXUxQKY3Z3cY++3JUGy2w0OW3qs77OkO7T3orwB0S1kpaIe21TeYBUnpBBt
8r2KmB8W15KLtBmcLfPoFsNwsYDqF6FJdyDVctkj9LhOl2mRWOPlegxTH36BbnfE
D5ozcWPrLz1PZQOIe8AaILS8BZLkWZhwMcRMvBB8X/wTdayYrekF02lCEHYmSBQS
O5pQKKOXxqxWwadWnLouremO2t0not5aFxtI7sVANNHCz5+a60cYu6g3Ep0ox6u2
7vXsLjSUOUoRZyYvCyQ4BPmrtb3oHHWLIL/VF3xytsS5Avx24dYvuJjlm/5hvGwu
4+KQ1S1c3XsrQwsIPqB3bS4pQP6UJcH+oTl2vUJtIls0uF0+jOK3hawhkVQSrdT5
pEzsMLrKS56pknabg0qwEOM+62WMBgzaotqvsEa3aHCKdTKng4SrMoJfXw1ZiAEW
e7+Na5Yc9V1KXRnH3qow9pcd1ycWnVzEJXOKN0nGvAhEy7MeCP2F2Vqw67ftd2nq
+7rN5kQXF/XcPABgClysM/fiMJcysxMLZ6+sJLVOOTa3aR0sp5ben8D+LySnJqHt
It4VepaWobL3YRGxXXLsHj31Md4RGZdFTeGCGnsFDG7ujnzXlohWJNG6YzwgjPYJ
wFMo9fa+STA5B0280wbIxiZmK1QsSIRuhZNNk13E7nYp3pO5qLvmhngh2QpRXPiN
XlJ24dsFrJr+3IGpWSoLfVVzxfb3ZjsVEjsaYcKa3TSxz9xcWz983hFwk9+wn6/c
NziQOU8lzZhfHuQpx7a/s6ZuksLa2Xs+YNw3OySB49CFAOuQeLrL3VCzwFvtW3B+
fqI56nEADVJ1fle3ucCiJjk1mVT0YB5tl4knP/Rf1Cbsw7BEElUCgH9w4cxFnavi
Cd/hw7IrVhUnl9ju1PrrBzE4WFmtmOP6kwuD10ISpHc127qzRNoLrqy73xrELYA4
jsFE8tNaoeHwMAKhQ1W/hKhv4A46tNi0KUuy+E36rJntRkUr9k83xJvXPShjkRBj
F0n7U0As2XJZpeMtJoNg9A5I80rvZkCxOXcCWRdsKwEoW4VGYVAufLDB0U+XkB1L
WgSqbcf1POk85EZsONcqFj/RYJYknptQNuc7Z+lytOhNpgLdj2iPKzD8TxG45RFg
Uj5D+e8oM/VfPOx1lZ2ut9l2l2d/OglnKrNVzBhU0pqET+0ifvn0kMepCeWN5CGb
BMno5R9NOHp25ycXjSalrqM1QIYEBcXyGc7mI6hYvuAle1xz0OUgP8cQveelaUs3
jqclXybGohDAoseO9VyZionPvs1AcyTAskKKAOi8EFNwk+l7jOpsmMU05yQ2WrGZ
JDLTEh25GZKmZWGZe0Xeq2eq1l/EdpGW1APzVL9cOCG48DPbDaiPaf7MJ0/d03s9
6661XBIIjfK6bzQxIROIfhqnK4cCMNdXXN7rmF1UlgWHJ3Z4A1II30aXjTTqOvEq
FJ7CNxzVrynU5apdmaf+961q+U5fwTtOXoPy2V6/GsnU9fxgezGU4ADhypPe6T9U
SPBibMDgYNUrX86qzhdpSnuQ/dcJyxvNR5DPmpQi3dMV9YIgUVIvhsGFAJr6iC/C
lbL1WCO9olJzBdzT2KcRimhLCnL5Nu+pxoKmS9oGPtiSUpdVBiM01/fF8KVx05G8
trilRAjcP0V2O4j7ANqocHQzfLbC2VaUuFYagVBNCrcTO72M2wHUTIHrq7wXdqN0
UP5ub6f2kwxU+YIB+aJmc5wCLLzz3sH0OsrJoko0uW3T7p0wIdnpsMG/vYbcjWSI
WJybRS8XpH2mP4B9awYAansOa49aKdIsxTL0Cqdvf8vwEEK5OOV3LSRCYHTKIXEI
poHlZyjGdnuShRREkAN6Fat0pUUiUK2ApdJiVCnTvrJ+qND7CoLWQZpBOXaXzsYU
AzqehHOerHjohDE+D4Zj+koH4WWoUlGFKg4sNmBYOcNiNRaypntogPW+IXgLr6c5
fvLnYD37Mjw/KVrwvZfSkddCpveNQ70SyOpUmjkhMcUEqlIWROslPinoaQF7WZh5
/5tOhAkL+vLbiMFxH/xzDriwiU4eZqgesONl2I5bStOtjwmXoF2SjRN/jsLEejn7
F3jKJ95vPz6vyZSz20wZ4VuvvSZR1DXvTYKrHvQeQKDEPLIe/GgfpLe0FKmjtxD+
tOzDpJN1uTQITyIMfFQGQNUORuzVKi2CILXiUpZSxxXxGmyJghTHPwyex/HZ2cQv
xSLBMFw7TyjAdIc43ZJs6y/KSgeV0y6vQOprUgoGVqKfL1mVTcoS8+6O4aerMQy4
NyAG8Qk+j+LEs0rY1S+9hNlwbMs3NkhX36QqfRFt8KbLxY4itcnRSqcrRyNVTcen
BJaio7MQxmr/0usdpnaD4N4pxXn0WyHdAo6Rfo9F4bUQJoePUopDTUWymC50L1R5
Fl2HB2wks0S0AgEON9hGGQuvT41etPG8Xr+BNabUke2rTdSn4HoqoHtG0YBI2Bia
ywXEB2vzDfMYjYDvkUvEUSrYOADGti1R4p+bOmiIpQ2OR97EExWs7wEv09f5/ng6
keL9b66m7iIe8c3+Qz0P8XREvltdriuV30wyfJD8Z4QXP8B3k6tlvms7Nnmp0l0H
deFaBZT6x8xAA+5taSSpw8UCAHHpyqX6OhIFp84j8Opz5WfpkowyWCc0Jt5CfQ/h
G2PK1Ovd9iN3xKn2HUBIhVjBYUJXZR9fZcDh1oG4JorQxolxsUUBPyqUvhLHxujK
w21NIi+6oUUOfyoFu4f66Cj3Kduk1OWAPIKEgqM/jEkphQP1HkzFJe7hFiQtVNXU
OOosCUUUjm5mkeqs+kOMvomjd8ufZPbSF1GUhc0e96lukoftDGHfvnJ8BdkN6I34
8JOhHOivpHK4dHT3l9zJ1ZBjrLgF83QZSqX4PjABTOSeQtC1rUlcWD5mTWi3FMJl
wK19DQs6kaX90lCKtuit76FAgRnh3VDxdGL8haJnZHFtHhpaNulmzPxzTe8VcY1a
+oi9H2OXhOZlnuEts9U7RyIA5aeNd7npRuWYf4hleC1tIH74Fz3xDVmBBl4BgIDy
6uug8dVRfsFN3n4xNZAfAOaeHICxd/esraeSiTG94ElyUIYj71+Lte8llB2xYPBF
6mnC6+F97GaBEhtuDGzwUi7yUtb+sbDvWw3IBogSPt7JIJqUygZgK0AnWOgsXJB5
Desrb6zoF5Ngz1M1ySYU/2XRnRDGjvqpB/CL/ZZzI5scVBhVDPeiBdzgsYgHlSU9
8HEij1dMAPIaIogON1+3ESgODXnO8SeLqomhVGC9HysjA/mYbmil92vcKYk6IAA4
NklNPXPt78ZXswl7OyxBrV8XmHBa2drLz9Tx77nLqAo0w/+wLFylGuEr7UjVCHVZ
C5rnaD5k5NSL2BILVTnZJQR0HR05k/DGxjYCUjiwE8RN471rpijsj8oxnneSktvT
O6FOrtAaulu2I/bZyNIy5jYnNWLivo7XnKWDXLvGiDbWgd/5PD4BvhB54gPRMcDh
SYezxcsjEVUvXwjemXR+srIG9+0BBekqSjfnEQQKM6SySZlMXSE6iA+XHVXFovTB
+jV3DHFZtA5BBuK9Eqk0RH+dU96ze9SLY7a8WvymoW3ZZe706hB8A+U7ZAp7EMDv
svUmMn/Bo7AsEDxRCaBuA72dyDB/ZmlBJ3gj+PV/UZAmoj4IAKgnSNLAfUX5fN5P
qzIZNfWnvPMqWKdcOpH3tgYC1M4WpKwEkHavg/fi9Ur8nl+7PKRyZgOdYlStsNku
83eeCJpI8VbT75mpoWKHyt0+urqvSQXIWMhTKT1F9/0zgmH+fyvzA5o5HDwtL2A4
bDvDJH3l7Pmo7mXneR/ijAtCLvbCTRBbReOllcxxCUtTryGJY5zfDBiSlhnXjA2u
FP0CCzBsJIhIOu8ZjKX96Q7rtyhIkmw0PQNjIxGb+aIJkT80ZWvardyrC4vUR+Yl
Z4gAPLmEmLn5PcxDVipNmpU0gm7oiN4zy7+61xLfZOIHCTlvYhTwCdKHvifFWIJt
K0Rv5JSt5VpHsj8TWpjtVR6S1zfWPLlB43FvHdBwA5zFdaQHmQIFAgu9FiCgl0td
XUxdAIq24CidSLYHXbup6KCppo2vxdYCpf5IhQPY+hwOiIp7SA0nhF+1IheVrPel
zff3e/AXqXJ3Ec/6yNqGS1YBYhsUa3rZo/6btkTl8u33PbvUKT/7LiFWNp3xKs/t
zUhUGk7rnNATcitHrJ7T6DIFtEt6XfUJdI52Ko7UE0RXZleVLTVK98XPIUFW6cs0
PJIGdFrP7DYndoQ4pZYVU+7BZYvOdyig1is1JzRebyB8P3O3Bhl3u2FIO/7KapLV
oKqEq1K1aEaUa1+Z7gJ6wXIUbqhwklKee5LiBR+T31RTXKIvo5Uvqlx3LxV/yHEa
y8zBPRlyPt9N0CKcf31uRJqs8XMp+0D+CxzzZIzhYf9e+w/jP060mBPcc2ZIPPwY
ABNhevMgTvPc6FguALGWNCsG04qOk40uHy7Wo4sok9mJcg/4aJKkUnDRQMs5rEOG
UHoUolPvW5gpLvBfO3drMCI6yIXNNBh6o7TtIeXZ/nHWRub3m4yL1MCgNf3M5ZRv
zwESehi3XIVfdEZbV7zc+pIVH3QK7hF370vvxezI2l7uRD7KGGaFK9psGdKFJHab
gzlpspbN6eO60hrrde9a44Ai3Ik5eoJanrWUQHijR/cQnhnV3Ihi3UGHHHA2pX6n
04o9sYNbWP5sjfM+Kt4xAtwiq+t8wsQ/ybKqAhEnq4gKI7WanYyqyPFpj4Wg/DwI
hYcu83AWD0wTtyntkz27rGFu1e94ub9M+kywdB+NlcdDMwH2jSUVbJACOsJnyZqB
GNVrTG1YWq6TZWJtFfGsgZTOZIeXotBk+D2WzxJi1CP1eXFrh3/7ZvQE0RZ2Ei7Q
zaJKUNnTlDDwj5anx/aHTG4uX0xPh1Gmuwm6olE+lSzsuTz7w/RZBguSEyBe4476
gGGdi6WkppRXlMl0A/r2yPiQ5JCQYl7/VW81RQr+Ofs6RL9EjkiWoREzYV2yHQX2
MNMBadscWrs79IadX9mgXQqO9upv83pNX33Yw6InrlT0QLKu3phNL5HinFkM2k19
CBXeDxWQ3mCYx6Cr/xlE/4RM2qOW71J/dNm85jdeCCPkNwZRccJe63R/HBqAe9YU
u7GkNDOHEmub2D2AUVAmM/EfLkZ9D/aMy7/wfyNL36Ck1sq0G9yBmlQSi+1H5wbQ
QJnpGOi/DpDxk3jL9o7ReDBE+68282jNSnNhPivNCq1eSWVkR83bUIcPKfoI7nSC
chCI6zY21WCeQB/xuGs2I0Q8sLoXA3KPcRUaZU74Y2oBCO39YMU7Fvnhr505kCRd
/HocfSylxxwJwPL/M5Jg3ZfK3pfPjqzcSb9ylkx8cwmoguJuJwW9eA1TJ5PkfJ+b
9IPsd6IfbnPuh+sf+Y4+TqbFKEJxcHTKfSzghauOK7/Ga/34H63VkzXZmlQaEicF
qUC5ioAM3UR7/mWLSSO4KprmHHFwKOlNrxP+WAGYZkeE1GMBvqfeMXK3rLIFPgIM
F8IMAWxU0IoiImate0jzwRE8/GpDSzr2kCsAsWjplZ+OtaUHaxcwTNtIkjX42LX1
6cHKy3Q6/v5C7GThcnNX7a0+Oy+RMCwpzuNbhshPoj8uUWwVX23spPz4/SU5r9G7
jNwNlIcKwZpA9oKnU3e4O/e5as6vxD5zhKh8IgkKhZO0BMcGe67qOXkLrAhsbWtg
NVwaUTETkMUUqDXMs5ko2GlxcG52CosqOMg17cRb4JH4C8sJUGg/KxrIIGYGlfFd
fy2nv5C/048BRDHn88EK2Z9giGHDdMskV+TNb5Wnb0L1gntTLkw13X7ZH2WF6WWc
3HAEs83547647eE7Q2pLWhVhDrjryDf13HEM4HDQRY9HCV3SmHmS0Eou4tJ9FHvh
LD3wPlYGplbdgJVuRFL/obtAezVG1GVazYNRux9Y3i/eVryOvzDsJMR8tf2+5YmW
yGMpKBzrEuF0XelayBHtO2dEtHSsE8UVg0SOdMseBgiKBPg3J4jZBDN611N78DX8
sthnCPoTguesaW44FHTfkgge0SNG4BQ9wEyoZgzaa10RCzJ6n67F/baxo9IctCZ2
R4t/ul+Tb3goEnps54r5Q1BHTGFlT1xWNvaCk9LHu5iDLaK8gb0FmnmUP0ud22X7
WNQQ1VZn/iKeAl7kVd5YetaJAGjadB93MVaGMiqkrlEMcB3wUiwX3tUQMxQDepqe
h951i/joste7hfIRcLPoynUAJK0hQHrDcBavTnOrW4T/PVC/KciDll9bMikSAdoJ
R1xxU5WFGbIgTvCGKZxJtGxV0UY6pARE5MgBbQCTMHkTu3e/0J6Nr2lTcVcDQzN4
qO45R50gqohA/Ul4VUAK8bASZQ5id4ym4dhwTf1lDv+GHfkDyfebbA5g1ANbNsnt
68sXj+yANfW9HKxhq7L5+zupx4mSu/G0P/UXCLk8r78c4Jv+tCLcki0/kASYRwut
3KRpFu2nqESTx6Q18yvNi6WUy4KBG8TJRzaj0cpz58wuWolsF02TZcTn21KMxBH3
MEgEvpDimw/XZQQDHIJmaYfewjGhojxJ39WxJczlIabq9NpFWmPXMJrvGFYN3bgL
6yC5tagft27appggzjcVMpw3nPNio3gExzkBNxSWEW43D4EpkPgQU9TQwpNjmQD5
JM7uu5Qn8TC4HjusTuivSpsP+Dp6QrwxhDPuuE44WKxeu3rVE5ICZ3DoaMxL8lTc
CHRlUve81I1irFpi97vY0x5A2dFgrb86f7aQOTe/YGtsWFwuChy0hCVaDkZwbHGY
dHhu1bfACA6QBFjLj3nmKfwWrrmzk+da3DfZDYyAs00ZHCq5/H9aLau0hOqi91a2
LNGpNOtaFunjSF4gRSSUzHj5oCNMDhp/PbpgsebLsIg/JAUYPiFnjenHuFceJV2z
ReygvHTy2VgKjSQdlWC5nxKTGEkcRr6iqI3dbfLgvdgU5efy3PzG99rCdYeaCtnn
oOuZBqeVHfeL7UMYhv3ZzN3I6kfWBLUrap7zT/VLwAPoDY4lx8Up0x0epGhb9ehc
EPQ/Dn0s8YqNBb8VWB/6QykMDnoG1C9iG9ormaZLsHTguUPJK6tz8ALoRMYpBLXJ
MtHs6I2DN/F1KyAVAy6OXJ/hl9EbRq+uyEctwdDqTaeg/OzhzH7KhJ0i6oN2NNbM
DVDUTaa3mn5vPr6JLHMCG14NsopzTyby6p5kEbrPzMyh6jOzbHcCc4U8aSdBy8xo
cJGL0RVDsV8Sxc4ckTerV3IJjMrg+M/s5nFoVi94VWq5tu57zhTB3uSwaIM21Oak
GAxiyq9mgoFnmXSd9GXYqnk32Z74Z7KJ3ZTjHddNPBZV9SnRnFyzJssLIts/k4T0
whsJnJGtbLROV4uVvL0qIxMgTVi4f6kf/1eyM3MeN5uSEl7IEfviUivt9c13e2nP
KqngbsDcu9Sh61QIuR8xrsEnimD52G1Tj9BSndG5k4qEmM5fn+YMsduhZuBtTA3j
Y2Jfgg7LDh4T95X1sBBx5kP0w3lEOGtnHzQObpj38BnhOHswMXaQsCPtqYRkD5L7
5iXKdu9pQqUjvcaHknWN/luVWGEjgsrBif5XjoYPaHC6nGDuxUZqU7v7hV9wBANe
5mHMk4i9r+H9jp03b9StHQ1+FevRm6EwIqvGkknZwXZhGxpFIvbKr026BUsoHilu
9oHNN/jJYkFf/OIPX2dqhUd2wRltJP2zCEc/fqfq7ILA8ik1NZ3xa9AueY1W0J68
XOf3VEVm29/FfHdFBol8gqOy/hsubhYBqJLFjpshusyXI+Zgtk/TiD8CwK/HdJm5
2yeKM9zaWnmJToqijqniCMT/FFaczSkmK7tFwKGOxRz6AhwKeR1y3M/hPxiUjH+H
CLd5Wl+PfYpbQjKiLM3dheML95P5p3D4KqA+KU9nhbJ6a3GI8SsB4nzJGdh5yADd
XqJ16zpxHQwpeVaGmGLqT4pRx5LaHlhAxt7K0V8KV9q9vBZrbSDatzX3+IDknwfd
Xqlep61f3Zqt1bImwxdrJ1486dL02JRmIVgZm/if+Ybbwt9sgqUDAr7+zPyEO9DS
AIJrHuUDFyAT6EO21Iw/jUc6ixm26fTKFVY9Nuqk7oJ1caNBu+HAWnwklEIktWnS
BBFs8x1OrAlG6qAbtxiUtDQWzz1DamzTgfvw7rF4NU2EjbQXf4jkm1FxyEyEw+o2
SPJLcoU/QEZ5wXsqI6D20iFxeaSffSyHyJ7goFc0GELYWYlhb/0JTjjEuda+bzng
1comalMJaM2IEnx6PWvyEgMc3ZsWJHxi7FYGgp3rS6c6skAELesdRTvzyn7s7MdI
fpCMHRYVBQycdxOe4939dbjYTajr5eCFAkJO89PtS2fCmxQSSHDMtlbqKBfE/Gnz
1VHpGhx85hkWSw4blLouw1zc9O04qx5SjevwHUTsSB6D83Gf724O94RZrfCLYwhQ
BLznvzg3q4wDcgVtVw3jnHuuD6wugAv62Bqob1gOJGlGqNyETLYGy6td2GJvvFoK
2JWktXLr8Xja2iuU5mzRuHIlxCgWBMPfwujbC0fFs04NlKPhoEMMU+hFq8R9YxWr
ebGmMovZwwACLpFIqhn2offW0y6B7bRy4J8g7x9Oc9UVRcYNGD3wHDpk1/+eGZOE
v00vSQFrlMmGsXOLgpVuS0vH+qMIPCYhUObGNRnqaG+4h2DqVVZS3nmDUO1Q7t40
hfKmH/rmxJUu6VcyMGe+Ri0zCKOReYhCHO8sK25gM0vuuqPTHRf75jHMmbpU/4QJ
tTr+18YEuEg7SzrLXf3zBZBXunbB99nIKuWSaSfvvj2mEiGcC9iI951LS9+x3Fs7
gTQ1bCIxVZxMci2wAKtIoTUtEWLIExzTrULUX2h5WUMtmQjjv3ZgLGaKy7+pOm20
ftgfDtDAC0gxF0SnCnYi/tmcs+meChAiUa2MnyxJ+FPycsDObuueL90jMs3vZJ3Y
4T7EJ+OJZqpBdoPHTPi2aUWbYb4bErrImWIh9xc2wqKwu253eNqcMDlJ03SiX87Q
9CRlqbeiGNFq2y658ikMcOhBMgeER3diToh0Cg+BxWYWHHJXb6BB2w8WydJM7hRe
SS4djhiHQn7GykyJKt9KvYUt787S6E5iOUFAHgUXJZeQbgWc1dk7fQalQfNrZm1u
yFUflNmchlfOMbsDyDs0CFPW4l0683QdMjbDmrruBDPHZmLWe0LS/vvofFKIeyJh
eCsSiBt/aB2u7AWP4cHv+EogMMXHBJlZTug/sZ6I4zkRmmKYcf/WU7JpAU7F2cjZ
/pGJCOi3LsONcg32h7Mszdix71B+NuzMOszSDvKXl+FVTGiGgyB+FmQJtXg+IqZk
UHsjl8cKrw49B0aULaEHTv82pDUS5cB4GJ5MTNNcrHH2EDWeLd2+DXPm/Xr+ju2W
zKWyPCXIZQ0ITkSGB59eZZvEhDPuTi0YGF4+n8LwTO4Z1PaYSMX9M8l0BgqNqPia
0ZF/Z1W9m1MTr4qYjvbF48O4scRZvcoyLT8OtDBQviVoAba0JNShOOe0KHDdEIy6
MgVC+h//ZWT2CoIuQHblzAFeGLfdVaJBq3TjTuWZzSPi/7FqgkhNmr8KfeSF1USm
7xDKJwumLV6ltOo5BMRKl016Qo/bAwCqYvuV/Pub0RRLmxdrhYvigTIPmE6IaEfJ
nanauZx06n0pJqLcODAnKtqEAvjpkoGPmatBDyTu+aqP6nk8HmlV4asdul+5IbZv
r66I/z44FU7qlJxL7tBVTSWgaUrUMLfM4ra3fVaO/4qPnMldjrQCjdGdCQidZD4T
RDFQEGOUTJ2UFlMJxa/JSwlWdUSQxD7N7qoAufVaZM7ksRHC3quzsWRZs8SMVLDK
6xhcTiaPAQJvsMzPJcuCP8W96P5cFh+eKDVMA5KuqV0gOQqQhP7KBjX0XLy3EWzt
Fv7ORIDKPZe2/ywmyiSqB6sPKUHSWndPASglnUwvmhIVxOhZidMvZuJynq6KddBw
GN6/sGrhJ5k7ue93BSJSy0CUeWhBXXs0RnoPqVY4fHODy3zP8o62GphQxaUUOsHD
mv/QpqcVC+qb6CaykWsYpuAF7nviGvfeAHsiUDzVglwPSTGqGP9BdYsVZrYYmLBn
CEOh7JzziSnwHNPylLCRsUCe02Lpp3zzvgRt93KjUTatLZaVtA0J1fN7EZqaa2Gi
43Y7agCpaKuEfPi4BXHamFF9jN5wh6c2JyKHZu7Wc8z2Nbluk3cXHCWOLgZ/+TEp
HCvYcFND8zTjc6+LjUQULlOPNpJt6scb1Lrkq14t25GH2WqUv6YTqLRvaPO2dFsp
GE7cyJ+G3ur1W039ZeAcLkfsrpvLq/QeF1pKI2ZS1wZZmqX9uNOgFm8B3mKQS5M+
Agbo2Y4irqkIUKan9/YFJUgwtj+6oL+KV629vcASJInS0MZmWgJrvglXQOuwavzI
ZGpdYhtLnOdWU8Y9z8k4A/0P9r0tBLNr55r9Ag6n7/szItI6MHQR7Ng8kGsFYoKM
BfIMUpcHl02x+42ae9jSPLAcOdnUFeY7J+6bn5FZNSL3meDKVTuKPElDpFuixYsC
ybNmHStqR8+wfopCjYl11CuxJ7Sz2N8IRfT797+yl/iEBBSKShIvUfXjSpRY/ncH
rP1d/fJi0HvNljlneE+lghcuG03o5vZz00X0M3zcGbO8Hk4Mol+SxSqQyJbeR22f
vEC/nkKt3rRszty3kcpisujxirSP2rVbtlWtzp9s1S9UWVZxnWVZPTwIAAdXvpxF
T40E/PA4NIBTWoqqVKoGmRna8icTl028nD4XNK/Qp1XDkGpKeI7HywEAkGUUnuP8
4ri6N/Wl+yFw3Wrk4cN6SZTTG9IOY7ohBn5J3gDmh3drPU8MxXHE+4BUWDJQgjgY
DKY5j8+9lUQ5nFd+gH9J9n9SCDMwRBiT+m4AnZhh7d3HxmXKjb7aPrSERISha2d4
7mMBLtHwDSq+ZacSyjYfBurtiaTwv2fTgsv1xcpoNKExcvfslj0PEBV3sze7lh0a
q3njTElAv30+e7PaAlXK71ecE/29HeiMoiVRd3BwHrkgd6tu2MBc36p8xVgOQLKQ
JKllT1KdMyFPbLfupuJhbx2ExREiWduo1pfX5ucAgY/Su2Oau7OMAPtneaoegNoJ
I08I98qkROnetHi/vlq+LvNWn1kwKqzXctyoh4jIKUmIvrO2Q6KXC0AQkKgab0PO
/l+P9UQKfYMh0JS8SrKUZNCzq904WHHN2wkJ3fKAZPbpMov3idasZLZzyo/lFUTA
BKNYbG9PbzHh4JtHJrbTqfWZVh8wedjpT8by5aOPJ3QMjdRtO+AGgwrr5maicrHY
51/zlU2gQH1pqVkZO8zs12vwTT6W6WctLCjBv94+Mr4fwp636r668gQGnflcGrLF
kruFmwixKOHLsY/MO71j14NAUeXE0BJDLRL83SD43cnyu9huqB10MAGaBWT1ST+4
/+rRsxetJs4uOdwSJ4826G908bIvQbac+aTQMmAwOKrrftAqpXi21Et5ggql7Oan
lFPQH9Jn0wZ5rLEim3TukmOl2Rdr0Fjm0zbWEe68FF844FgkmuO0bhz2YeM24go8
caTKMmFzjoMuni0AjqABBEbIpjdUgqj5gZY4EffiO46zxa0Dk7ipXa1pybmTW95+
luwcR7Efkn8uEGvktDPbs35UBGtrcRX7FcBvhfRuJj9cjoswetorY1ffLjQBudQd
d3XvS6J+tF/h6btrWyIJr5Zlq4TCk9Dhj6wHSCir709vnvgFHmg2xNLtw6O1r/Ox
+ry/rEv5rAxf3YvswcUlOpof6Lc4/vslbF8kg9v8+58bSeLtwmNUwepmEYXATh/B
GR72dMLoC3knkw9laOpVzTB1lAekrly1PIbIltXecHPECb0R9yv25F+9h9++zq4A
h+MTBz6eoWZUmieuTWmHF7y7KFl37b+Jl/YPtGopgdeS/wjnAV+j8zoFE33fxxdj
Ztny6hefPGAh7TwD7zellUSDV01di3/umldwJOzBKERU7Up5P8k0mVxModq753kF
/BfbnwncVFbA2URizbOjwkRafJA+c2HzHS7EISDYXPLlKYUTOiuoUz6s/3sC3G9R
86T6H0qBOLd0uxb+apIfT69Ho+Et1LDalya5c5qlsdjweR7jpo9xtDeG76LYVZkv
kg87Fz4w+kuCWnNEg5ePuANpVedQOFMgFyjVDjgHa3P4fqYICG3+hMh7u8uI0Zt7
sndsG222qxp+dbpfbJaaaiy9aP31Jn+UI3mJIhjetXW14NPawoLFs0uEKxebWSnv
nUlbEEd6QCVF9rv1+Zk2bmVjAZeaK+oWIU2uvIVuR2TJHIXYUi54bU3WnmbECPPz
g+B9DZhvfA0zjRn4UhnNLwrlstlJbjk9znGATbp6T0SzC9ckD8rx5JNJNTEymAZ1
YBHfGyeB24ri7j01V0M1FcnXJ49IA0de5Wp925FCzDB69OnQ+r5uwNcSs4kA7PYO
bKP/TGMHLhg9JLctQ4PY9q6jI1zYJhrfEbEuKyL8g8D4lWQQYj8apkH43dNhxJ+L
QK5z1DFtspNIrGLkcGEChh5ZwksbOz/5fuEKjgVAAg1Gjlcf/Y8ALnbmnG/x7LOG
1URJvzO5IYcD+jGwUroZC3kk7pVuaVqIO6DO3cEDfX7kB6l67VNFU0JikCJzeH7A
Jd8UZs2iZcLM/XgxE3EjH8Ue3QO7ghtO2FbF0NMgPMCmAqhgXxdyH/1KMtH1LUg6
9gBGqh9DHZZ1HjgRb96MKMla5hpejW9WUVsa8fja6a+wjeQVjXW8oqcmche2fsXj
jWTCvSOAzgOwHVJs2GeWt4jRHZUYAb1pZD2aD7Zce/Gg+R8AZSSu8OJ5TQEPkrUH
A5uMmpXmPeqEyOl7wbrF/8KNZuYS/PmUOKgDVVQ29p5eBj65K+BGLkRjqjlmtmTp
Y5x0QyD3POdKAJu5r3zls6L9seT9TgCNEVB46y0aTYkSV/bMTECs6PX5Tb95ncok
7/k1L4CbP3kguF/8MRWvsS+Bj8uA2ADPZ0FlaafGwpVTRMBeBQR507d59nN3oqLN
7waFZmlPS4AnHeeYj2R7KCYX0Jt+ktz67lmSE8uNwrtVgTG30D3u+Q+a0h7qDtHA
sDL+ua+X3lO0dCUQOBGR8MhpK9d/NJ5LqKLPCxLTi81CmlaE2xvsijQhrBoSG1GE
dMjEu6tmy1PRgIjQiNWTAucj1fDFW3mdl21kJ0FKXPvQ+YvqA7T54PwQonLEUbAQ
7LP53WgaCEFoBJ52y9BKwy2jf+j0r95VpPC0tTLsCvDay2Xu72KA9LO31h7nNZe4
KEgoH0lkOkc6sv/kPjpf0djdGYKoD6fGMv+lbfbpcWOJiQ3adOCbTnhJYbEGFet7
rR2sZVsDebn7AFF2eGY//WvN9zSADBsLUy70z+wntB6FQ8OoVQ2+umFkNklEAv8I
0EZkbvw3a+NGIvpXpOBaQ8Uep9WDkPpfWvJVVNmYMP88G6vW51zQOlxV0KtgZewU
JhLAaKQroCPO3Weg+IrSVhcVl4ItQt5Vt5T3Zvy9BPAp9VymUrzJOA61HgKCu+oW
ttM5Pf1hlKKICEoesRc5cBmasPuylrazcoEMkJsb+r1ET9xu0Gdi+d/PCIaMKb9y
m4yw7tIc08++zA7tJLZde3/pinthYoxTUnFJuYJ0H7PLXA53yA44Sg4UJpyWfKtn
xBzm3jgx8NT7JMUBgT9Ijn7BueQS0nOj8S9QX/YIP0cYi4AQAtKCcdhIBlXOZwIL
g+jXndlZbHAUDESv6lMew2mUuzG5qfdpyKeBjQz/olkDCRYi/Rj5CZooBxMNyZmE
d5DMYPZz1LODLy4Bo3DliZfwg5CbvqqCxDLbSBLLFQ3R08Y7i3zhRXoMQ6d4VFDO
JhZzBWqRqOapAnfwpG+vxmXi9dsMYSrEgagqjyQtCfFVxJK9pUcoIdeAaBI7qJXk
A/xmZ93WUiVP5eC/Lt3QTyJ8DfDCFqk4x1EbBdZOAbmE+pxaCI6LXyAdB4uIaRhs
6WXpTWVz7MsDZ2sK0muE14PyZr4Q8COavl+8kPPio3VSLxCnEj1qzMJ+AoArm4Wq
OcONMdxhPmrZ95/lfKxw1IKFUvjNp7P/PIdsLq5bEZTfOtY5EiZxpLqHqcalr9s1
I1f3O2DaZCtdmGIq42j0qp7uAWutLPUiNIxkCboa+jorwQ/rWpuOuJFBvP0qPWkr
vwtHhtgGk/Zp9gtyf7TOwwYzOmbVQtMlm+2+14oO69qVRR+DoONinO9czynTIIsU
9DnKAuOUicvaarABG61i3NQCiVD1LDwKyx1JdQgTC4We57KxUEDm7+z6uoSp53zr
5TtZiTeuaiJsXvD73q7RaXFQF8FHHNXzsmSBlsjzi5sUxe8a7egZlQWxFpj4vjBe
X0jeoo/Iu0ICXcJeX1xT2Oyo8qHn6dckwTHfY1qldoEtC+CQJ4LTen3Mao77A7cj
LD/br8LqB3VzC3IiAZdEJuABrGUpA4ZwPggWv+DbWcYm9lLZ47BsbAGYaZYsSOkI
GJo5albQxP7j1r2ccMxNTfRgRLJlx2zmxHTlqT/iWrWEALaMDDeUfuo07De3HWpd
OPcexu1h5q1tTzsN3irEUk4CdJjNcUWt4LDZuyK9VpzGGxQhp3eQMzJHTNejD69T
d3RD/RBidZD7RltYnWRaMZbAytD7TVNxvUbmTYyqOAhTMmvmjShMmfEO84ifQfuP
WqqhvXS5dU3V1SYGEIhdKTxc1m6R7uOFsR1YMhDs9dyfropAS8m3jEYkDh5wYbFP
MKJBiQqyamRV61kWfo+VGstaYbMKwcyxBe9+tpVZeG/3iYBgLyIlkM2bC/YgFMRR
yC2hrI0k2DjP1/fATTfcUsk6hNREUaSaSfDiMe3gN6r2rlXnpDk7cKorTISmflGX
cQQjXf2JZvi+Y5wYpP1u4xANExbl3DUystCL7vdNEscKEI5IwFepK/82bqzp1W0O
uatc/WSS9bWLQFa7pttidpIQiQ6f6q7p3PDdiMrM/nSuANyn1ttcWexxAM9pGpwZ
rVXPhLQ3o/7UuY993kMnJAqUcfvCN32ugyN2s8aZBUcygFGIgRSkmWQmtZYNowsH
Bxkr9WUF4XcatEZsEpInvn+1clVPKLmzD9grYW8h/W80OtE7Tx9q0BgbZILP2Tvr
gs7ZcyA9MO3f3udAxcqeXlPH/oAXn4qHUF+B0f8S98Q3nM3E+PEnUHLu1rwzIaGI
iVZ/qXqB6MVnQgVuViZ7eJuDiI+ZMXlPsxtXg7Lr4+VjGQ3IVVfhCgJ35WiIUKKm
EvyLkvlT+33Ql11V+K5U+fWCa6eWbXIzOzw+BlDEJV+dBeYkpYvAh26WThFyDi6d
QVNimHVpdXgCpn0PnITJ5Yzjgc1J5MYJIyFTLEbUsJmY69sHnnl2VryfykZ3smuX
++NjaEAW5NOgKIqeVh5tPomlFR8zhBjn9Q6Ofoz06zzxMlM+2zkCO07Mc2ATb3Nw
iHgtgdAMdYAcJqa/fu0jiha7gnXf4RR69px4sRxkQpG1VCYgsEBnz6gTDe5AMoVS
n/lohFm+JzkzAidgsUjMJqw+LRdU8tnJD6MGlagXjxICi3QKlq05wag6eo0wJidq
n6hvCihiNtujRqBuT13YwhHuBP8Th9okz9Jy779HBzJsaag9n3/EKVCs6AlKnHJG
dGgMmQvEVSOdDNlcItYkHTC7F54/izEWzwBV2TOCNwvM5OutAapvic/bbVSOschn
V68n+GVaVnSvKkZIaBtjL2x/0CWZMyToaFKzWdviq+l3Dg0XTLyjvt66YVnNBFnp
xS3169I+icnSzJ8JgcidYqCIncmeE5JzCyFnIQxuqHrH8ys8FHhh+MFSy1xJguqz
Uojb3FT5ik9AMbkcZqavb9I77tCK2su3qkoJnQeSVLq088e1eHbALLljTBzl+PQz
nsLtjgYiXrbFs4HG8fkj8fMMd/9jKXp3hWiipmBVAHqmdA2bp8k+Y27iRq1vry6b
4cNpKz9jcPSWCiIsGGsV5S48jUkXqhkbRNzA/B95+Q4dsKbftOThzBOt5sS+/bFU
/ZWXWPgINlebGYrixfS9XEXcgtnSqxDsV5M7+17B5BeTW9s8MtKH3PODVTYqneLO
Grox6GxQIEABRWiWCZvfiWxFemF82cVec6p3qqlBtErPZVMpgRexnLpXG3ibB1Jm
r0FKzR2NVZ7dg8paHr+g029IHE12mWU8qmbLfXeawmO7RUmdSF80fCEd17A3aceI
tbaWCqYpG9tZWPt2H9H/TwJ1jcGGwmSAzCPmzPeuJhDhnxr0M/muyLCisMYQXkEj
bvbepCwq5uD8M7qv+iXrLFzMWz//p7SPpUziH/8JgjTXP1pvXdeQAZd2Fe0IOB39
4mD59nDRhHWBumw4Pxqb5VeNY+7G+7wW5ULsYKDf49Ywl5xgAof3upYP4keR2FkU
rCwGXjm4Qdz+IwwYoCtbgfH3rANikjMxc/cBlE66GeghKzluuw8UhdmgCnGDpqTv
jq79AdNaCbsG4663t3YIat9cQlhZRfkN7U+DZzogDdXBrfKcNm0kPwujULvQMuVF
fExtImGyF5iVxMZiFkL7Nya2fCGeUUCU+BNhaXbozxsZFc2ZCbTlnT7sCcfzS8lz
D0kmx6XBkkDwkWyraJJpzzGTz25VI5WImcxLomBzbpKuLITDcHNz6VpbvcyrCZRZ
kxUm6WG3G2Lcwm9a4pfgg/PZY49kPoKAan9KYM/aOBc2t1rep9mtuxvTsC5y4LvJ
bFLC9dwSyAoGkKP9uxdrELS9pID9Et0zE1NWdDW834bW0j+/VsKCb2ivkfS9OFls
Id9XCrZy5bgwg6UkgOYkt8axUOfRhGLeIgPHSahZvP91ykFO8Yn/4Pu7TFK/b9rH
7m6+exZjSIQgxlOeLhStgmJZw6CdFbb0FSMrUN6UTHBMsQguBsh2i0XWcPlGe1z5
i9TsEdlJJgR+Juc/dYFVQ5vQhEJB2+xiZJjqWoDlykC459K5AAwvlfjKj8kryjb0
Zl9CNpz2mlsGVg60LkOKcgpk+sxM5XMg15bz0+vhDRCntoIKaGO2ALaUmoV4Rph2
pl9oVDcJbNve7a800eZBrIFmZWHFb6/AhosemSOnS68lZIzMmZqqDB/e2EtegXBq
phdfYBio2HZXrbKwlwgLN4n8qUFtnsIahoB5nvTjVwArATFMHfr4hPRLHWGmRwPv
FD+o/pEKg0wrKIRE0jQ+F1rjpPK1szOqdWQSYRT/HAGzT1pkMQ+A+9mlxE0t2Ajo
QNQkT9GwaD30La1NLCEcUAgbT5hin7l83+f2FkMemaM6pYaQq/3yYNB8bctEUmnj
F1Cx9dVOmLTyOapIc9NU4b8/K0EzUBl8LkzXE5DiPjgJ33Mu/bTqCzl+AOO9OiGT
+WB8kKVhlCKjY3ssT0rCqIHKzvyd7l4EI67ethWdXFhux3cE5o2m9VVWgh1apdD0
o3CFGbUx4jCW8hwKMxt5TFn2a/4ceDeziINohyDVi2LwpKmeshgQ1WFvDtumzMFJ
bDQYSnkfKGeYbtYvlbrF5HajvCuPz8UbgJIsyXti9BstJZglBrNiBRgP2T9Lp2Ow
kO1SuYMvJjU8XY03PwRnuj8dXrtZWvOwy0Nu5qYx32zw7KvEtZgaGpLCS5b+ykKN
x27+d8bESdMcSqnE3LjgSd8WcFYuW6SuV9fMHZhFe75lreL74DNN8xJwm4HFHQTz
kg5ErPkpwGTnDLTEVwjxheTV1Q2F6i4AYiuPQ11Y6SyEB+IJ3tJahXwthL27Itgv
LvJhm8GNCjlhnu6vCbSvL0J4dg4Rz6QY4vu19K9Ijv7CaV8o+dIrh/hOwAjI1ta9
nCfasGaJ2Pt3dD+jXWhx2SQOSlVavXygfCf4FGu7vgqD3HG54cQ0aaWQjUwBnqLs
6KeAUAwMubMxJxYo0kRcTl4ZmQEYWTtiqMZUPygBxqUxq5pLqq3+sGFqkFqNLl6u
wBik7NE/iHnIxW2rKA0GyFqbJKPEc7SGZGt+aNFFMhZPVhWwLXP2k9YidXuZKmpg
5Psz3cSeICtYh/x6+KosPyzyIqMzxm/4ZQE7AXgczRBzdmjJGdvLDr6HqxmX1/Jl
lTfRXc80bM8dYqNbzbKOKQDUx4RPJu03Bzc4YKR3tE8ZZDKpQJqfpBekHOmAYdGZ
yyhfo/TWn0LFwlTCQ4+SOsasFkJQ97ce6ez7dL2ER9cpPOctOllZpAJSbgQdfteH
M7cTarNUwCdcMm0XxKWnQVe64+XdQxR19RAAC2tVflaiH2k4pL/1qEKly3E+dxGy
WJrRn5MNK4iLi/Xk6GyfV2HF4rOP4XioN8MIqxXGhV1Sr4KpjqNbjB4fLUcxu+t+
+0a2hkFjtmz3vwdXF9kaBhY7hNMwHyo13r9e14eRklBJouJvQ38l4S/lBAxbni6y
Djqo6nVFlLxLP4xK568KjooOdkY/WExEf4JPhoKyu/lgY3S8rPnQTWP4TmG8vGoA
4d0fOlIRNTZpOMER3U9+jGSlSIc6ZsbxdLg4Z3c4N4HSw21DYzzLFeg4LNMpxCo8
EeEnmHy/bjmdWLRIZ7HNvdXHm5/XoR/oXUP0jarNPAICNYT/hYlwi+0IPwS9g20Y
F+i4a2zdScDN9YITLVH4YORJwcMM50OXChtfNcpzYKFKxCvX3ST04vECSUXJPFkv
iwSHowJ1g6z1ucEsiO0w7YSGJVA1ofF1delCEkVWZXepGeEiWKYabfyj3l26jV8v
btZLrGsy0qfvGwu2k+sJQsR2rX7vwofG742GOV8YjhV4PQ9i2jFxZ3LcKCjDu9cu
TZ7IdJfmsAE6JPEkfwOLlk4gx7qaKRmJeI/KPIz+YKT0J0u777OfzL/kkVNeQAl7
uUc1pFki4VTRsGkzMED7kaVP4/nlY0XsAPE3ax+wesOxpVnpNScuyKNKVQIjavww
eLebDvnvJoD+7iR3SMXuou68m1F4K+fH1a8E+unowA6QnkBY/9EDZuMFsH72YZKz
P6WI9MNovUNs3Ul1fGzCtiM/4hEFXQhoyGTld3O1eqoTt9Vjmgr/B6QsmgTL98sy
l3xyrtxB5bHM7jj4oR1OJ8ZRBuk6dzLYhTu1Szy/pEDcqY/ep8Cc89oy7WyA7BGa
3so3YnMJXUCS3KQOMJPbk82ok3+O3tadnvCexoIgti0y3fO2JVN2mgUxcPf4x8rv
9HzKrZ1QJk56H5jonwaqksMzLRGGWYN4YyFWBZwpMi5sBGyaUH09deiOS2BnYRec
bZglPbsItguNItUI8PI6mGfrEig0bxB7wRUzPHWQAb9YH2C5TVKw/qDoaIsiGt4v
QVK62VIk8kplK5ynV8K+VMpvQk7BvQ+KkI0ra5SrhJWfjSxme/h+FXpKnwd3jGmv
0tzRXX6O0oZWpuSKGIXN405GaQH4N2Y9w3dKXdIzmY1hwfTw78FQqaUMJim5Pj6t
m2qCsMFZfrnJs+CtJyQKmhT2q6n1yEEWnyAWOz89JJI+ZRbotrvgEOQpIExBKiu3
zT++t5+Bb53jfW1r53+NSs23z6db8U6/rDTWxJWkYmJa9emVfMtMJgi6OzKDrdyg
x8G6ofR/a/AAAw/vSiTAj4eg/BiAYsq7vD1OKxRbB9XPWed4YfuOcckc93l76rpp
qBsd9qc97fDMhFCj8dDbYBn+hVAQYsVMIRWmvJ6XE9qVhv2h8CfigUD17kXsulOE
9ymmcPHiS6JefbjFbe9SHMhgvvk9DHBSHmiM6PyzA0gu+rZnjSFBE6LbONM+On0i
3n0CsRufQDaX0KifRo1Dr37P0X1mJLttyo9PrV9rGm3Aa9AacyADeF5cAXR7oFwV
LPbZ2YlX6mqXKr8cbSQpOcUkhzTYw3DuElLS/x5mdjPqgKC7CBM5NWHBh8g4r6su
nnX8SdgQHBx0zvc7ee9nGO39cWJgsKBm2kuffHO5KokU8DRuuoUkD7ExQQgDEIvg
PN8tx3LpCFJJvaRAMU811Vv6/bQ/Z1uXlQtpuFFlR9OTm8Q7SYjB9fbUjSCvk9pv
ZIxJV60ONMbm3fSC2hU0c0T1gmhJWb8iZBP4u8wSh8OhhVIUC/YS9WmCkqa6De3g
Bmk9jvTfNKKp42C/mlytJGN33duBBX7zhBUYBQAB9FSXodGin2pVXXxQ0xOf5H/j
pnGD4020LZ9+DpKEQbnO0PGZ0YDkmnrW96XAdpiOL63Lvep4TLNdvPXasHC59+eb
PRVjs0x0EupY4m6NNUE09UwSHTSlTy/MvPVsI0ZAF1iHRrhE1GVN+CovANAWKSx9
k4KEYM0KwGrqkXQMhmnb54Ys4awnsTZHSR8C/cKS+Kl+5b1c3Vm0zZ38tQ3OXlXH
WY97WKsM0LS6+l3IhqQGGZM/EKlp6FyAT2oSZUdjlonAoY3F4wsIZ8KCPfeP0iFi
ZF6ABULWX3gomEIISv0GVQfSwODSZS2S5uu/GWKwzb5W+tpw5BnATAbPlXHMSlcF
wSXrwBDqfb9nzWxkBz3Hm1bHuACyZaHHXLh0Ob1yr2ppfwMaQ9868RsjGu3QXewU
hUeiYcJulaUf/b3M1GGVVBYmzz3smj9XIw4NxlSXHQd4dczA2MVltqZEWHtBHAAd
EiOJWx3SUSh/Yi3lPRBR7jKdw72cB14EtICBTgbgTflR/deNBlqmPPSgyyvwao18
VOOyiPoAz1glllBxborp/Fg21SYYXrJfwpbqn1b/Meuz/aFNsAVbxiyxoEb8f/6G
8VIFPdYJkTW3BSDorE53iUc9W5iPJl5psFwk4WCSYJM0S93Iw4bFrPWAnsXsTCYM
G8bLcJnx/1QFOi+uBcKSM58UoVgUAI3MkCK8hUPAHzXp1FkS4DaLyPyRmGz2jbMD
vllvi0MAyl2o+7Pw3WlWaVPt/EpagcReltkKDVqEBEMhUzu/r2PXlh6Txj713Bo/
an46Evl3OIQ+Ps7xuzn8pGjMGINBvb9UQwDOgv72oelJDDN91ZGpsb9wK59m8s9n
O2haBDoiH9yLlf0s3E9Lw2SGrDt3xEoZJEyMr1/XbhIcC04cTYPAd4Fih1hZ+MPX
Ky72fzo8nDSQQW82OdR41kL9A0hVywzvjVkqzpSQIB/pfZIeClayp0L+n8gOmXFn
71WeLNxWmBsSVqNjrnPJZ4jZVYR/GSJF0fKMUWooTGsM/+aT2X4DfNIQK4KwlCVI
1m+W0diIZ0+uTXg8fXWdVXBZ12FfaXtNMq4NQW5E1QntboApJz6+dmJwL/BXugn7
t7rJWPnnFhg9WO6E0nPDzaReyOmg1ZHSJtvwhYxqA9LcDy8fC4FEwB+Evj+d2OyM
Ky89HZc2AYYASrF8JRfDFn3W5S+ptwGzX7YkbxeofkyKv/HOQUUOoNQWNjtNvnrd
7TYUtfLw/yFC9/b4MpTnOcoLcndnTiH3+uZdY2HUnbgkRn3/8sPlDp1tU4Odcn6H
I2TIbmPo0j0e4XdCaalhI49A8hwYZDcYSX6+OlKzdkqlAUAJ8diOUKQCrbPLTokD
U5lpWSpsn5TJUitWGn84wXu3MdnW0mRUcNi1TE8IKgU3IYIaJlKpg6t/lT/DCMSe
8hgZfu7LdE0vEXM0OjyJpx8UCt/anGBa4cL/JnXMpT5fU0KO/6zFrcvMv5o7dCqC
hCTqwWVrpc/JluIDIG1atLZG7sXE4FHC7VR7oEMgkukuhhNb7AAL+HEPzyLDXL7E
2+hhjf9/kBU7vpMv90NwQsgvKQUzxShoXZBZ/f/1C1C9pB5ly5wQlmNfsQDCcDl1
t7c/QCxkWdxaO5drw4xmfPCIB8hI/lLg9AaWkpOhyCy6LSe+B20SHURCVEa50XPL
nTi1ptA7C7JePacFCSS+YykniwSYn086LUossV8O+hH/9ffk2mc3MKyE/yNIDKpk
YrPQyJ6WhKE5KRkKRZShP716D4sJTR3QNNTZ9xymg22aSVH66M9DnhAhf511ClIr
Pl+7GCPU86OzWkJLShYtvXKqZmy159+XEgunx90h1Rvu0MY6fzXZ8VkK8yQLpJ9u
O4u+6SOjlKAjCozV7LmkPhPVQdMjkXSUT3Zoxv7VkTrCkunWJZA2JZMVCBJ42sDR
rRNiKCJc2SYqa8TOcgj1GCAEh2yEGmhLq+woyS0qbl36cxLYXeC9oBrhvLR/6hdU
Y5HJjgjFUJDHBBHLAtZWnMoGCRGxa0hw4lh9URe0ki7bZ9Lz4F//jYjHru4WBQFs
yn+QuZgOmwfL+499qR64PVFIu9r6MoMoUyvrCdmNY0jah7YmH5+//vXw9XKlwDe9
iT+xzQCIrhwffzWXxAhPX9H7tiZ/HApEbknnsynDA3gfG/DScLKCSLj7zerKKL60
UNzts2HL5lT6V4104S+inxZec8Q3ZlPB3YjxBdOHEVKXqD44phQ4jPwC1gf7d8hz
u3OTjwfCmOPQteU/3YIBOrVgLBXPwagA3nT1TjNju1gWtc3oomgigddMkJZ3d5Vf
nuriAoVSVmP9pYxxOwQlWX2sFWFo+Z9vX1jSo6DT9et+aE1PTOdyfevHhcyVfwAP
+0tVzMQlAd9L8hmMU7X0R9R482/1/W8r2lGFXAv86s8+P4pmIC71G/UNFIKOc6Jn
r3JQfIAgUqACiE/J1pq/QaP+T/25rezS7tVDEnjNx2kpCcTVwGXEm6ald/QNG6nj
Cdj+MZwetpNdXeSmnByCxGrhEaz0tU2yRGeaN0urHHCb3IsB1+/NsNLnv+zGNMgV
e5EEKsKpKevMxF0b9c3yHgWa+UQKa3LQ+e8DuBbJLdELFoSSUja+RzzijsZJ4mT1
hzQFABh+YX0HdaLA/VblpXg4aSGjiP5l/n04PjQzaeqww4TnhATohMm+R3hA9fk4
x8c5ER9FY0CioeiLHad5cY840F6EnL2Tcp4Y1UiYG7y1S0OJmLESI7mjjHo77WD/
o3Y8uPucCpIvEvOkT3plEEu3a4uj56lVva5p5Rs7vrQDctYamLOl1ur0rk5sfJjx
42vZA7vM2JuJw1IHQjwITM8pcQqYp64TtOy3m+NJw6xoOif/j6cGmhspU7ukTnvY
CLb69Kdp8h3z0T2dcFiAIrVQ4j2ohvkOfyY2n62EfRbrmLr72mBloetjpfNCE/kh
o5/5ZE5n51fxCZveG0UB9ZRLzlh4XvyTOevqwBRSnPAE/1Hd0rd+QCZ+cJheupir
JraGo46rQ/vFrG8K8fNUZYguwDtG1y45USI+aliqVLQfxN57zWwANLQzdjwberzD
gzISYofp933VbzkzCrpC1R7uBRw58nrP1PUnA72P28UUui5w5UGSpdo+VpJ1pOGk
OCrQB49o/VnB0y0zmLO2p1XJRKIzVSynfBnqduE+UYpPlVrEfgn6aPzFnJuhH9HE
04tUp+MoxpXezhhb+1zruQKGXJL2dNw4o7Tr8fcCDANFs0FVbJzQNpCd5+Xr0z9b
WRxIi9zSSkzFp19sGm9ZXTXEB9BsZhk7rf0jcHTSRzyBB41ViRwhPJqnxUO1SVw2
0m6C2jBheVqF7w5K7IePlj2tL99tInhNepm9qSBGZsLUPH7rTigCvOm8Qgwhleom
eizNavjkiJQXHzqLGLlsRu0iBNJHZBDY32CJ8yphAfq9HVkHvbiSg8UvCq3gVMvA
r3TsjYKTxsWC98mkbM3a9GvsHwr5mdM7lpHcDEzgQbNt+f+TZ/PJgOfVMExw+UTB
WboAYD+D9RM89GXlMLyWAlddVwU57dhhPSxmuAn2dUSkmI468oNGzaa6lYR4cbCe
84xZBx3WM458d+9jYnCNYRKs0A7dtdl4Pf1AdW1OmPJ22pny1cRqZ7OPyledG6PG
QrPU0C6y6wqHD0X3cGGgTriWk4tvsw2tKBQw3GMmSfVRP4EA3PaxHOCwPhL9gdTm
zoizCAoFyQF3hjz7EZKwgnbJ5HLHCZVXoZidoi0y/7NGYhB1aNjePdi2bxV/pZA9
oNA9s83kv6KPqQDdezFjg+nZqrbW08EhjKp7jzBcTlEEA4ICEj7CUpQjU2z7gAVo
Op/0X9A1I+N4MHXy0pS0CGg8fKhgSrw+P940rAcP2N96JPRbRWrn93/ZUdXAtbrF
AmVnLpSuUqrgxbyKi2cTGyKNZ6rmO4ErO7LpF4C/FUE4whWqPv7gNtt7jsRwlcP5
KYsqDKjrDpvgt+cKV7dT4WTBQJBREHlIuoNfgSBY6qXdoK7ZdZMEeg6FqTWVheYt
UQ8wQ6T78QJmgpO/p0SoyZodLgVg6WcBIC7eG6sDV/hRhr+C7eVBZ1ReRuXg4mNv
JRT7Ffz4H98OklzNXWYYnJ5nJOFP/pGTraQHq4fHHjSClylTbtukKhu1NjGK3ZlI
pLJ2n+BEAWn0es62BFMA30B3tlKxtS3BI0e/hXCcrT1I5ruTip7jzt3XDSfMa8ED
2SHL3xfoRn62nlEz6bIpqGdhRzJj/COU+qZ1QjdBYrFQlMdcqdJ/3HU+AbBQGPII
f09L1Y6p+l7lQFtbTOsjzIxpga5XM0UW9aS8fb0UazX7xJ3Jf9YQdW8MkDVDb0cI
5U5LEuq4fg71w6Z1enx+5kQRrjH6f9MeAFGUQ702WQPVDOd0OUGrCEYOZY4U3ClA
4hhWwBxLwZecvJ2xVcbSpWzhTSrhWbjXI6S+la1l4XjxK7GKz61KR5tnBvHoXTWB
8J6QQMxJq+1lgOzqoaIhRUyyoHFSY2lypO4ECNho/uLwd0zmysN18u4ccsawxmy/
ypjbqx9/QFFQdhiISx9WTbr+F2x5MJB7BHaZy5tEjRZr1SOTnEghvVvOpWPxn4DJ
/T3gkHsN9ZUzksZzeqdvUGXlwmDgwTPsHPBjQqqNSqKazVFiTZ0PmMQ6vXS7HSd1
tiyQIH49a4s/zQ3dpZ6cPRj3daoFGf2YVNJI4UlEQlG6yoYG+Tp1hPMJ3CCy4n9W
p6BfLRBt+DkiqnkP3pTfXivS26Yygp84RsEICBdZLpQH0Xchm7iXbs59b6waWVfS
Y7Ky8yz4Cezlq9q1Zh7liRUgK6kWoAcTfw6gGjxwonK9zOEDTaohl1ED71PUNgw9
t/Olk1PdWQV3LqL1Pg1gv/5ZxLPp+7t5Vzjv7LhjFUJXVX1EddE0AhInYjF3lBoE
GORxAiiS0rHk3wRJ5qtGmdGeSG9ybMf9aRDlsYK5iSt1c4RjFmLjekUxtOv0KhxO
FDpFYElCC6M6Hij7LYkatLPBWW/EiKhKGbIQzjGn2PGDsrDfRaVm5ig8LgQeu+ct
72AbYJoKhfwroKwDsRaoyhTWrNxvN1fz8lkq5nW7bunm4bTVzNr9+4riNU5+/i/C
Ee6YO5q1D1VoLYRobBS6VtNTl2uwdrdhslFVdfWqeJqGOF2qzSyxbt1UQDXjdmKW
lavkNwtoTM80J1FhTZemy1ap+wtPcQ1xt+TGCQkbJT3ipX/VyT8csJOBBNHCej3n
rXiE6Wz0mkJpwDw0oRGvPDlHMlp/cmRqiobWc/4wGRijmZVHy1Hfd+BDCAiUTe6v
fAJAsxMfx6l6fEQBM4Wwyi+K5twERePZ1cIZeFmPuBvCpkELB6uOUJj7j/6yE/ws
rR/5+gcL7q+3ycUlavXtm6mWexWhnCknPf15fhUD/vNWnJXd8pTB58k4P7yV3M2M
67loXgzxKxcEPAKZc7BNmCLA3BuLPAIjDICiZ8sj9J4rc4TUUxMoMa1PWtWoMzFr
7qxwuq85HTp/Sh112xyRyRjRN5OCn4Su0PAfX4r5j4p8bDqU0Gl+CUB5ypiekdqR
uAQVpn7DrvXoF0zYn+2KDKd+6H04g/l+oIsEqVYX/Z/kX0kJkHhNB1sSyxPlh+YR
VPHW4JMJVT64u1r7aIRB06VtLsnSVhAqSwaj4nX1C42oZ6bMKXvQ8uXCzgKQrqE7
/nYeP3L0UVFBbYzQmy+dMz1tYC4tV7FnkGxrulYg9iCDWXmC8/QLGB/Paxhaj9C6
q2R0fCNtwjUkepEfwS4ulj4umDj++bFK03Nf1dQl6uMLdiidD9vtPCIEUZ/HmOf6
mpHSBuKiqwAIonuRet5kMf9TLEn+PfFizNmmLNzCROc5jT1SQz8Vt34hx6d+1hdq
x9lxM4NkS1L45wstE3ZtCTgMvqxEvuQyZL6Q6hh1ffncouq7ZA4OMZjobq4UF1Qv
bOozIQgLuqZnDmVDlT9qrj8j2bPXwPCJooKlP+9ftGWslzUNJGoP49lf7A2HJ4t8
7eRs+1PwO5gs48GqezVo0tmAIYLnH6aIjukWTTctXKRvNI5VymREmVFMSCQcN2m6
ZUkQ5W5h9mQI5u+4U7rVrk6sKRAeeLFkNGSu85AQKle4YZmdaD1mEyBq91vUOhIX
w/OqK+WrfPyH0waxWHJhQW52rF7ddAvnGCm4q4gSy0WQMw+8VW+2FzCfoCtdPGpL
gMi1Rv3Evv+mhOI6K7T6QJ6sRNi1vZRNZetjq6A+rW/sSIFk1HJmh4zIxirwRaQ3
tWmGhJY2X7NfOZQlQRNgzmc4mgmrLMvUBxjvvVr5Mi8GiDtbnjP4a2N5h5+vAbBf
jt4ajhkpXkgazQ2FKfXPjNR0f4rehnNkJY+qOYNO1DJaE27fmqMl4ocws1En9rPd
q/ekMDDIMd56ckSo2bJbZMX8IZ/L1pyyILsLZJ8VrfkUdkJ5NU6WYBlskWdERI4c
P6OHJwUv5e+/wrMTepft8iiN9FAt5OrLCk8l/P6rD9bBJOmWihL0FFOKgxWW0Z0R
rVz64eHQt5YumQ6t3fvhToM9qOD6v/c8HFkmc+tPDD00e0jdE24OoVzWlbAPG2J2
21HUSI/RmluH8X6ccdiFmv3lEs7MW3BsdAEjgKGjUNeLpXfx7l9ADO9w0yuRlsb2
lU6cTgh62Qh9vHRQAdIGSm/tCJLhbLTbIYsacYELnt1/Q4QCZttNojpEN50QP46b
GQCJsxkT11eHFZ+oc5vsrjEkmoLUVwRWM2qTCVZi6dJxPTI2r1suPxSY0EE+7oP1
BAVcFOMJ3LMX7fhV7Ajm9c10yyoxmKIWxvC1Nq95XuzGx2eE7h4evOg+Wf6flPWp
xuWwlyBbQcQtGMjHYfFkbHdDRGMacovGw3cHAhjvHeKtm8q+0t1rI80oIb4ztJ/a
k7udb7Bngf0f4pUYCxbfPNuKaXlj3baQL7uF5xKltfuHQEb364V+qFAb3P4hRjE8
Q/lLc+rk6/Q5RbnwG51CxKf6395HuT5+sHEIck0SBCJr0ZI0Re366wZ1CwZP+wJB
LUs/7wXXMyAkl1kh+PGTKJIvmYzJoSU8+B1js6xVHS3T2AoLu35y3lzq8SdnggP3
6UE/goAw3AwdVQlQ3G6OUPobdxomcghepDIjaDi1zhdKjD0UeI0Si5jpS42qWvk8
vRhn8JkCWJCNLcFlViw6LGc/re/DmT7IDD2RmdGsflOPO89e6mt91euz9LdgWC5u
ftGxixP7bAN3BAQ8p5i6cWP9baE7ct52GCoS1S0iEORie9qUxqdCEi9lm+MXD8Ak
nEFTLWOrofLh5UrVOxWtQyrNOWYjQT9aih1yRWt/dCQJ/BoNTWuNpGmUmqBqV8Ch
veT0dZrOPYL54dmkF2TnbjWBYc6mAOTuwMY8yVu0YiyMcje+u+3Axqox2IENXYK4
yz5uupY+2gYST2gjfUrZDrsWq4DlsJBSDway/Pi1oTFpkYYdQMij91g8yNS2VUKt
wysU7WB0RBoa4Ts5VfATaA3dYEgkp6Ec7wfoqnQtgy9XOBPMaVRo+eABENTF4Om5
X3HJbZfRrN7BROAmLPiCsQuI8RTyybVAKT2IJGnDuKCtkK+JoLQnUQS9pfuR+ifw
YXEkSytmIxPKOu73BPqWkCRzKU/r2Qg2nJLjRj6/y3ZQhKCB+l1j/Zg5yNK2VQJ6
tesc8Q1FJovoClWuLp+txNmuFmZ+13K3UHBWo7tZ9vLSVIEy2oiTnhuDYQz+jybZ
9BPCVCyVw5f0LYWNwXgeCJKuqkObKCZ0esm+mobKq0T4WgOBEJ+/XPJJHsVZaCtp
SlCvcwLU1C0blBZ23NaoVBivrUWClTgvHaNnEUtDQ9vcbmkAQjRoOR6euIUA8vpK
RkNPLwa8S5u78oFC8vmv9ZXsWEcngdZ4v+crXVpic5uR86IwhGTuR6BlrlcXj7jP
Bw04GIs0CvdXpHuInbZFuAfxGL6FvkzuaEYNkg36afJXcu3WHtFGDdDqIg/BRBc/
I62ZDzZl87kewuyPoAmyFPJzEDQjC4Q0p3VwH+/Axv8yOeXSYN1ERYDV2hghDDLn
AZVn705XYbE17lyxm52ZIjITU0UeqcwnlHeqD72T9sGmjKGg+9x9fCfGNlL/o1JJ
oP9d8yji+0TrQ0gYqguqPzlkjqysJfnNSDmGv3Zs/TTGHg+Gsq22pP6W5Bg+J+HS
prSRVjxIkOtTwiHfUseQSgItsGqhorNEPtMpziheMrvMC1mw/e0uBGcw3B/BjoV9
N5dWG7/RhMLDywKmUj7C0csuNBzR2gKFmZ7zrPKqjAnz/T/i9pU248D9FJ1PWQnJ
KJDnmYIuNYE9dVFeDb107DgtvaQ32RYQTPH1leehEQGVoWe3yna96kA2VNBb4Qvf
BlwAuRIcflPNJAuzs6ezFIHs7lmPaxqYN7Uo0a0KqlJLuOT6GcQSJIB++09ZBO16
UM1PtbzreU0eFXo8YZPIK/B7re9WC1v1N4FueZxJjbPZopE8zuMlaFXl4SziwkSl
DX5dZU9mjuEmgDnBJxPqwel6+XYwpDOsfhPFGiA1V4w7g2Y+MvBrwTmY+SJBjdDk
P/LxPmERB6U0ugQuwoIBrfn1vYIwXSXNJzjxa6q6nRoYsWgm3frnxqKuDNMFX24n
vkBy7vMNt/73taq4PbP5ZCmdZbJMIbuk3UwpzJPNYEaG2BLV0GvMxBEtz2JKN3K/
OzJD+8ZMsMr7IDYP2D4JCu2IitapBrzyz2v1vcVOTm8xg1UK+uULAP1SlfkPcy0Q
K2uPBywH+MOBhmidl+dMD8rSDIlVMxfIqO4irgbHAN01r3F+zqHw7beDbGWyxyMx
3arGudFfKFaSRVcMkO4CHn4SHtmlLF9+FZQIE9mqWf8hSal2kpgNDsWjKbkvO/mw
tVagBHju1+eK2PYEBpXkUOBy+apEJpAG0emYXscbGaWItJUol5ShNTHVkOsWXnG/
PjE2AxRVleVl8GT4iBrke5KJgG3I/18r84r2hcX7zJuGCR7FFfvLKxJFT4nqTq+f
i8EDDZzNGlfLWbX9GHMpEqrMxaKxjqA9//d1i/B96GlndFE6W/y1GzZuygbGCKj/
/2neppK1qp5YHvfxM1xUxCgvHbOPVpQPEEbzYvqLs2OwN2CwYnifWow7YueZKiEw
pPXFA+epxHI/6R7xV5A1Gopm3mGr+l2zanf/TQ5nv3FHDMDzM5bOnE7EA7yJ6tzK
5a9nUPRmm5yDNNpACRPuJ4+OepAp+cBxPgYR5csRG+R/7uKjMWmid6RTp1Uus+NT
jKxOZtdZE4eq96AymAX+0laOwNN+K+S4SmAOGnNhLX8yo/oZ3f764DxZ3/qN5J4q
AK7EABaxz29BJPuYcn9cDBYqrqT4jHt9MbDZmJEoqsYMAAByF+4+aHXuSMLBrBoz
GiV4RMFW3sxXEkIijyHPKQLA/zXJQ8oRJFrjd0C+9nG55Cg+NYQMRkNnKwHnNYN8
3JxwzLZf82iYgTt1lU5vWhCbQGspxvIU2SWK2ZbBugunC9V1bIhRkLA/eAYTX9QL
8P2N0diZ6BA2rvL5xCxSSTeqPNgy6oigDjqHu/BWnDxuuUztocfMO0S144IoJYMS
s0KnrhHDEQC4DWmvgKp+KENOFgLnL4Yc/MGaRIk17Z5v5YO40wrJ9geyw8cUXztF
eWCLa78qu9ruU0jvTO7FTBUl50o5c0ylRRsCxdT5xPD38pBevRpiYGOEHRkVG4us
nznoKO5dqfpTqtlmyiEtBd9ITlnXb4n6XleztjQ2AxCRVSkdt8jREysCrM5rUpVQ
0X/zN+T0fVTKy1CW5S8xv+3AEXh7sEwyyfxZd8EXm5B+D+jJ6zeMRbVCqV2M4EPu
weDgYfZBzn5Sya7CY9VLJnQcyQ6smIHUT+wumIK/AfqX0iMcv5miamNo1Oe6bcBJ
QOvqB9DJke3ycqqeVEDwacEt4EHg1VXh1p2Nm1Iha+G1COcGqndhlGjn3yf8jHQV
QNGa3vVCJRax5UFJPg47Iz2uD2LyZVWY4Xj8QsMyWzUvtVC09eLkk0NBptfJzjnt
LNi08H+NmS3oPy2TlbVZ8hBhis12B4EppRXcS0m3R7j3GkYgV1zFHu7V0WmtWTvh
meDV0/5Y22JIKrfXCgURo6P7ID8TxYO7ITB1fPBt6zDp9mU9qgavYELoElsySDPv
R66sTgvyjVb//MZnDUAkWxOUqoHAFxdM6BeexlP4HRRFFWr5GIp8ALJLFcsdO86Y
9OA+oAcGEF07buyNiGCa+2hgw5d/PGLoYhukt8/X1AW+Aq0L6utBe7IKtW3trsuj
qtQIR8WmAbx3VzSQDte5F89PxR5Vs1PSrdIImLAnOi8Spjhr2HEeXnBr8oGKIxLW
ba4VxefUz+NVB4kAs+B+0l7dszX+VUjiId15Wq1h/7eeDl0a7OatNjgxc5Vn+unj
Qc+xkkTx/N205Itp4pn5WNQvax8HgYEZz2tpO/+2egpa6eE7XJUUNMxBcwlnBEVI
yanIYCiahNxe983FpLxQg0DWept21vWDj1flrOseb/d1p4IXXevkyjIZGUXL1qgt
qH2uImMuWeuP4Teqo/T4j0zdhsNmss77vmkVvHohSRoZH+p/t1K+l48QAaQ3RJkd
NlOJuxsn0yab1W1DzppTtlFku2ecN3YBEGGubw79jdfOIcLqDdbapQqNWXN7SImt
i6OrFXkZJMPydPVc0C3Q6SMs0JVmfEFQwFvjMGoFWinu8bpyLPD2GyP4pFHtVrw6
di9Tty6un8DXO+gS3gOxiKsN3L1VbEnERyyCp9k36hUX1ovh1nFxdfKqUa5h+AS1
wK8r5Hft8nJ1ZZMoXS7+OWgDTnus5aVRgGlZowiFl5es8RnaC8A9IOChJ8uSuFay
gsTgHKg5ieJz/8O1UVQCNuB4ChOgs458s6USVGjHMsts4527eEEDwpNzTgnf2LEI
L458aELaDUPRCZ8HNVuFpvdnwrFJsPRF8qnRPpq1QRja7ipW5F3yM3Jc7cf5qIDM
U3mLxlkUg1zRDzvkB2OLsgEOOa1pltg9nXWFgAMX5e+LvManuMOzPMDvul28QcQp
pEyBwgzqw0ZB+7epf78ZPHS/hvkBYzXWSK//bd8bY8WgYOKrPVXAYr6HjfjB3zR1
TAbNisU8bpes6Esc36optvtMtKNVd08FwDtBMT4wz5vGH/eZvHwF7QIBU6WWIThV
8VwHe6gMntBKfDEmNnhWiKerTEqhPiHqeK1MphFmB5WHcs4sXY596ps3NuvNh8sM
4E783I/Q6pQ8AJaKIN84y4bglkpugvmozWpgKOJ7Nyun27GVI9Nxfix/8QxPrczo
RFhfvew+GcakJ/mWZXsvQTZB0BxlsCNmPlpdQoj7aKgUsNJ9+K3VtHR3aw6XRWDg
CsMtLRk+gxMg0IDx4mjlIlfBqs82Wy6yWkjUuHxB+PPJ7xuTPJAu2V3BPjutT7gg
nHRPhy6v2qLVGyz7LFD68VY+oLd4o3C75wWt6C7cVTfHSbUE+rY/OjpwpNJq2JYf
WQ9gFXSpF1gAu01nxsJPJnl5dN7ehI0Tf5zAVMx5LYN4j9m/l2UAjWIUZ9IbHiRJ
xeyxHPq5wugkmN10oDhgsygalBW7y4TX9JKWzv8N6ow8vzT+01UTQ0uls4KEBqn+
4d2xQsfmfIfqK/stBRlCf9ykxdGKLT+waIka1t5ejI+PzIuiKcSYJIsMTN0DeRem
std0Xo8AHELFkGfiZGFMt2p4iwIU05hDEWJ+LaY9qJddRXYRLWoHiulqV1XkkeYo
5YkJVVepk8CVhF0FZI7aYR+XuMU74RbcceIdEMe7W+319d+nAX3VBn+oA7gAO4ka
uh+0/kobi4K414kasc4WziqYwOr1X2n7o69PtKXKOeWRq1laJehr2gQehjgsKHMv
rcBc3f+FVReuofTslH7TUaBDuF6wu3qSDpl7wJ3ZLcsAo3B/kU8HxX0EX4FiqtLe
W/zm7BzM/601NaZVn4WvJZ2OtIdry2NFWhgd+k3Ht6RS5Z45UOtq3mctqIdYL63V
iB1OT7cnYl55RAM+Uzb1K7n4RhabtucK2Olfcgn30BjlkAsRu6+YzA7S8FSUiGef
Sqoq57zW/ua6AlDK0oizGa7eJH7OL++bfchy/iAN8y8bXR/rZ/Jd2uiuoG2FXPF7
95+WEWcE9+P1ePaBD+ibKhyYAxcEEGOggsuzR+FzOJUR+5cZfoFa5duNhJCNVSLw
IJzTX2TUM01IzPoAkJMNk5E8TJ8Zl+bq0kEh3jO4c6qjhdFFhKSb3fBc8jIlo+CA
ic5g1wMtqRbWsSmLV4FoYVXdafanfCqj+VkJVW+sPXlqSmn5qt+t/HM6yq67HMTT
C/QuX4fWiz0n80ZQCbwURy3zKnhh/7SreQMDTS9BBGIgAXrktl1YimAtLbHpyXrR
uQZCLcC0Gl763Bmd80ylurOZccruGxgPXIi9nWb8KZC0nD0v+AngH6E+jbV16f8K
BG64SgxHQ8SAoebZPjsAORiW1ylEuoUmV1jhL0hNn2N94SMY7RRdckKxx0rb09j/
RzuQATUTo3CY1q/HaBHALTFu1XWESvO7hpoZ872Sxxv6SlYQr6nGM4sDQmJ7c3aV
u39uxULgSTxyrOV+3ZEcr62MrZeMFa28mj0iujwugy+IBY08xIZwWzEzu+kPjBTi
4gHlUU9RWJSTfDApnhTkIJYO0K75V4LyUkjCRvyQ0FSduEJ7s+j7/HKRHeq6BReF
4HWMasq0LT/muvV6R6cFW01GrvdSBU1c1S5QtCdFG4F+Y8JXr8wfUp/0U/tb0i1J
CYkQECZMOO51oi+wbVDFGKiEZ+92bykIOUrB+/aVY4YKknbLOS0yeKWjRSVQuFHD
52lXEKwz3nzbeBZXtmkAUq33wL7QLadG1wJGZqaKoJyQELhPhNRvpYBSFoysYTJi
AAihCTScJEn9zq2ZX9LBHdICHniKKioTfmPg1dLk8pOeZcVYgCNOG+NkHNnQXH6C
9J4U9sUq/3BFGwgrmOTDXlyQ1x82PI1IDO5XSroqx80RAJtWT+uprRz91j6NOlAx
bFWTyCHOAPAWzK3I4gdyLMhK8xVh4jxGr8gAGwYCcl1wUNWJIvxH+ORsmIXn+R81
sUdmFPugDNk8Ju0fsnYj0iirwY0y0EPovjo8Syoev3HrNSsAIA7uVXer4GZvI4Ad
tU3QMqjAEuooaLoFLKXsxT5Eu1AzKwgdOTXZNIRJ12YLNk56MVy6LiiTfksZTWur
zqS6fQhJgoemhRcBscI20Sn6IxA601vFSyBRSvyjQ6aE08gbbsNvvmnZm//eHIQi
exC/H+zU9wbtYRB7IAD1gmE/IZq6PlO8Ux3MixkRDwuB6N4lW2KNNQr4RptBQ5CH
hjmMajfZyvYh/iRrndoRs/rM6ZBqkkzNw5FotH9mcysoEm18r5AKp8cLissGRAQx
//RoOhlFFAtPaPUttRtKRTZhrgwX/hawgtrMihaX4wQaPeIBFfhK0tomBaE/rE+Y
faWzSrr24tZGJcuK7R1KY7sqJ0VE5a2Mu984UqOqWRVq+pzCC/WGJSXbO659Va4S
58h+eKRO0rTp8BaOUSBjFdKgGfqxBRfVQjLZLzUXgSjVthhUBdSZPAy5h6+C2d45
vQIv3Xo+eOciMmzNxp/Cd2LmJAEcH1W6BWJZI37yZ3QRSJAScKLy2wAOpTQDwEB8
PI4COzOv/W0ZuvTzJkOzXcr6qH434yiQ1SmxsciIWtPrLIreSr4YQA9sQseIZi9r
uy9SGf1Vc26wHd+DzRchVT10I0LzWbSWPHo3ycY/Ov+0ons7n2ncrpWwsz4GWiE0
YsyrP71jm8Mb6FghRvxv7VUisXSNEpDsPxOs4Or7zZL1ELsbl4yen4sdyz0PDihw
FJxSk1hp3rQ5sp7GUG3GIlAvb+nx5WAS3pUW0iZzIEfjPCkIDapqUtjiaZQVsxyd
3p/SLlUQXud7qBLczoU3Vtp71NVELA2ApVU0N+BehyFr2OMXr0sHjVGjfxTAgv8+
+7TfqGiH00av0D9Tghd5szNiYTDQN6MzhyKQpgY9jSVMfq0J1490dRPF6xcuOUzM
U4kAyA0bEiIrM3RVXoa5upgu05c5bMRbeqAglSR1+5rSj8fJepvRxy8tlrJYczc+
TumuFMuK/6G0MSGFOv6buJiBIA+cCsGIt75dkWOI4lhaL2Xz5S3UInpr5pEAOg0V
Nz0B2aQcJSHSn+7BynLkrtvFb8RoIRRukNe10p2BwVqmRzckM4GdCudTzG1n2tIR
IiG40s9CM9ur/+K3H9+sQ2NJ7stgZgCLQyDkPb97mEfF8LCnciCwSFedp8I2COEk
PuAh48D8Ay5Y1hAGgjwsWKUUwrI/PlXlToVTmteZTIlYwMt+LnZ5BkYIOmR2hRIQ
HEQrpxid1zVo6eQJv0k53i5zUB5YJr+Nh3zVb7C03jmO5NjYo9mBd8bf5lTPKpDq
zHIzlxacZ/coOY7CEjHXJ1CgUtlZWDZsFKVapqE5nEicLChPdiI75rM8yndBcS6E
/XXOzel8ml/4PQGHy/MKDV5OC/JDSSTwKBV2WfJjL3TFouR7axcPmXwSVv0KO2oN
+gIWWTL6ROqEPvZtdh6JE3Mi8+r9S33y+e3uMdf0p94VPQdNcKOns4T5JKW/j26W
aHCWuZcnjx/D9NQw1GHrsX3NWmAjfnfx5xqUqLza/ctwR4oC7k7W/yF5VI1W+Eu0
94rsIRXbT3fci9x7czP69Mf2T9QSyK2rev5m9kPtIM+N8D6TUNIDRLku4rC1giwf
qTVIgUpePdjfuVoc3zvWDOOjZouEmm7A9JEdOB7dn8cuIN7KGAB6kfpHn9/PTuDS
urSMGhdRjc1sRjlVDES3CbT1IbwqXYwNGs+lXt9INYG+iOp6oW2Sji4rstjDvOeM
wDJkA9vqtYowAHfEwFlm9H42rEWx8TfBU0OySP7+mDi/U+XWsL17B4WMlal/QunY
WTbR7tV5AqvW1cjdd29zOBMBMpZyVfhd4oM0Etkb82WkyVL+At8vzzHttmxWUjfe
UipzEnDZigwkBc296/3HPUE+G5wlPlUZiRpnoPxWC9Fokpzd20pTb4NrLidvbv+j
wjmqvsriyIcH561ACrV3spPrVCTXxqOxZJ8L8Lj3/Hoa5xt8l1v+bJerU2rTRqLx
WyyLw8K2y3Ll0Zm3AdQjPFTVmenE6stkutiQGvxGIRM6KbXQ+h+ekBChutwr9rtD
TPpKIEE77nnARo6jxD/S9xIGTCE196Cn+W+CRurZmCZAcRRtNKgyvPwL+cfMWvLG
TZWC8gdTPpF16eszmtkeUiiOy8skhIEi530FxhyHUKw/eTJ9gQPC51lEdB+f+myb
j/go+bsA8KmyZ04xU3NoyaRVpwQNd4fz9lS66JCPp4RGZAzqkEyihC+LxEWkLEC7
+an/fqr6YyPNqhVUnM73WIeME5lCXxoYVql39sd8/9CTJPp1QXafTJpG1mEE1Gml
+rtoa6qQUTnKZx02cKWiMLxUwYrUg4P871nI9dOqzPhAtpLjj5YX7nXqss5RS3CW
jt8LoTYfy7K0e/W5LDzyz0jG+tcPDOZssT77DMT7NHFV4jLyRc8KswEDKHVzqMO4
/DxWCgQpGCQrc9/22syYoh+N1ngdxrexGjR3lRyoN4qvQpnWAq8slKBHG2e9wm/q
Gm/7966TNOy1feBq/uuhJk8bFCuciFxXv0J9R2GIQjTpXV191txkdVR2aMEMen5A
YK575QowUAW8yNL+JcauO6i9D87wQxURzqLR7K5ofyDw3X1l3aVfzIRFTtp6iJwA
5aq/r09hn7Gn0KMRiFJoSyNBmJI2/7erUZELGE9e9HCP05QifZIBaxwRKEmCYWP3
3oriFQKAeBtRm1S7cT/20/conieOJndj0VZz5Ft6LzwMvQqKJYxu9Oa6UCK9Q0nq
MgxPBVxJ+Mg7gfwqESUdQdeaYGYSNsx0PCmrRL3oLPU7JEm/LgiJwQUCHBhkPANH
ctZSRqVKiA5Esv36bG+QnAJgbhLQJ5SFa4EQmTaljUPrPN0gOpHpmcS0Q2+8Wv5u
0gSzNYGtvgJmFkeXy8PWIRsWHkrui9KceYjLVB/g4fAobEaCfdCmPP+LKilczOKS
BLHW2LxKX1EzMtpsg8wR811FPUWJOLvj2f5Es5o1rvPOxeYzH5sRyYAhdSvNYCkv
jmWgFKUnxKK6cT3CZyplLUNC0n3049NpMmsewXlMYbzJ0qyOl/8aeSMoTLlpBw4T
gVDGoDCO8TEnMIpl/N7MPwHL8zkydl9RIn/grVuP6y25XBlG3q+vnETV5Li52FVY
zNq4P4oQ3fudJD71ShhsppejSBkjUp8D05tcPv25IBfh8PVuEcNLXyeFjY/bAFuX
8t3ZBtqLlMyXIe+namEqFGpbGwnupWwdECFZOqxhhkaREOkwnA7QxI2E3UpWvBe8
EiL7DgZ2Q3O2ZtmH9WD30DRTyKTHjgASOMJaIORHJQEalINBpPZ5YvNpBxJcBji1
OYKNKMVQLw68wrc3GwIoD3oiNdSll0+NWvBJJU51msl0yt7K9IAeRJaRfOiZ7UBP
Rx6hojNMwLGZ9FnTG1EKZtUfW3ZO7UPBJktfzxrPRGk8wgjpO+i4uCL54Rorqst6
PhjGdSN860XWIvrViMJ5BM5kH+0yab/6whd2bFuoQZwctfSxOcoFOtTA71EwyMga
eAwh2HAdWrYJpcykhIFsdDoZcmDuZF8DltM4rEmdxUf3I9qc36VJ672O5Ba+dAcZ
Qz8D2n9lTiRcIdM5i6K0pjTKgdGUhsxt9yYhW0KByUvOHI413G+j8lvA5OghbBnj
FYbS9N91ISGsYLY5LC2rowieWwvExBlwC1dqUR9odWAmleKQnCBU1qhh2e4wRx0C
UmOWKhGRuUvSRiUtqeIRxiRUUw2nBuOuyug+DT6pff/le3xzBNcLa29ZPp82Tmuc
prHqFyNjyE2Qti486dprfpfK5hiaGtjl3tJ8aD5+7VsVrgMMjg1DwtPo+8GGMIvl
F9t1ln9gYeralsjWsbvGOogcBkDfzYpHkcYKnLgeJG4rR3/9dmAs+5WGhugzddHk
a0x+vW3IjDtlqadQempX0WWqz5fKCShgtcA81ml2BmJjog4wv0wQdbpcWiJvfesE
WbSAwfyjLUHA5dehdp/AmpNP06L8I9SaWJzJQtQfENf0jS794qvzoLukh7xl1jgt
eDMC9Ab02xbbvPFvl7wPefwKKTGUFTclM7mWxGDX0sG3BXFrL+oaPwxt6LS5QA+/
YmRgRHs2QjmkE+H2lV1gVRLvh+X99d/WL4Yk8DZHXOUDWc/bZvSjjcUHTgjw2y7+
k2hcIify+JTSR9pr5h2Rbwz4I947zRm+yfO3sZ2uMGJU80ynaqSEXQhPKYLCqiSB
9Nyi4ySLBf9SAT2CipSoVBQsjgiMW6/HG5tEeQsSDRbIs2x+MOqr6tTA47hC9PRS
P+PZOQLBMxyA7GU5/9SrW9V3zbpZY8v++8HsQs5sdFC1BX9/BXEybCLSTGwDJ8A/
DFuWQ/aeK4/I/HJ88R9Nr17NbUZw5LVIOgwCDONM6Dc4hs2cnh2Oa9/+d3mUXVts
r37fw0zq8sBfKpXgqKL2ISFtXG9C4paAEn+68NIwLGzxpexOpIlFwzuFzTzqPquW
D85JbenYtrtL6BE1U3eUOwuLc2XB3MM+Cl+hfXpGeUh+LqzjvZkeVfcTMGiaX+MK
+lVOtnKeAyovXevmaJpo+UYf+rey4kn5a+7ce1G3TPXZMX+S46Qfe1ivkVW9FfKG
5aaKoqN6MHK6V4J7J2TWaDjyiLim/KKDGZYI4Ej8xOivfda8qPR8Kos1FZJRLG9D
2FC3H99eaD3LjzFP82fDdD7H0VZo4MIFQ8f1skVP9SRHL9ubzF8deNn386rXihir
Y7FSph48YPtXJkD4vpqls9+JpkUXbl1mirdrpkOm5kbnKOB74yUz9/Y3PFneJUVa
UyXoIsgFRiQ2mFw6Py1/W/b9CRXKr1xMzZwfBH410LrmieURFLE0R5xqHjLFteYM
BFIZ6oZqHzwBGtSzWp5X593bEFeZA5aRelX3+p6PFg9qTb658eCuDIOrMm1XjIwx
+hZlJSaGQLe68dMj75daGBS9ZCl0os9bvPbXDhhIwilPdutHeeuDXKoZ4d2UfHge
685lfIVFt6EZV3Af4cYt7V3J19vRAK/jd13K/0DznjV0wBThgdQKMP3RbXCW/UTm
ZH0nmc1Sac0srN7DCPJIY3DO9rSzUfBdYq8Qlzu9yBRTv4PeZmgwPCOC6ZLbzmAF
6UCx114VFWI2ml7NTBVxwfCPb0MQgghjqBJJ5PrC5aC5e972SXzk2ETFDmUDkY5C
pbUOnmayeIQbGga7Z0YoM5GfCxqOBzxgAdpn+01G4FL6uNy9+1dTGZoKfbEtWUp7
BSsL+cYWKRGJCvKtNNAOclHDtgzcUXcB65ZQp2Ve0+yd1Bt33+heRQa7+wJRKMY+
GlPzy1nCOM4Uxvt8MmfvplS1Zln9zhRHs63g2yuRTH3Y2hQ05zzhR/Kobt//Zy6F
b5Kr9doo5xGed3OsTjHLH0V9EGndbpUmrc3tfScgmMgpyZFvEHrE6RYspZ4TkXwo
3iEogUdkiIKuEGBMe+Gdd3XCmL2zXbFaP5/3pgBuFUB+8A3xXA1yXkmkpH6OLLJr
3DeQMCygAqYxBqq1dby+DIFM0Ax2GlNsvA/yTbmqmtoXiHSkRN+89QvS2CJS16so
k8qAOMNul8k+G3dAEgIH28sjDfWQLmvqGH2ZhovLQceRABl/qKayuxGsqdysC008
p9zujeNkPO7saaVUM5LrMkM6u2bCUyaiWV0SpoF6EjiTHhej5x7qkhTOwQtxe89c
q++1H5QGp61Zeg5aqkqoGcaKD5nyKiG4X5hapXh4NTe1Mm/OR6sSLsAGF+rzKe4o
LCnAqJikqhY4KiverVwinp7XHUtx9vYnpTheONX1UHM3tKXFdXx9yEuwaHdCyVdG
xlXJMFaltwBZtLpc2HfYa9f028kccpY+F+2cZrq5GrVVEqG73IqbXdhW/CCDGIJ5
0tmzliEX4ADhj6+1DIGGrS044wvzjMOZNYpFM1mIphhNdimYrwuXG4Y1/jSONvP/
z8UttGQzg/PgZzYhe4ZVfz9SYx5s+VYBAcK7P2PNFT8DilRIjXouzubmoxEylJEw
NVW+0STWwFUHvnf+0Rz1IKy3Eg8doYVInAxzPiyyHpimTH7Db1xfVtD/XV69IaBo
ySPWxNOALuJojRfKAVUCd1kfzwQfA/EZDScHv5RJM8jqT+qDxrD9Zt5MIBH/zad9
WPs9oHeOJJ1SMo24j0teXxVPHjxoBBnx7VY/+pCy3rp/WHSZm8i6+IdqYh/gyeWy
RmD7PDXBV+T7+ou8e/CRV54O/srR6wloQeayrFmKfsl7lmhP7dE7C7g8HQWGG82O
BNW0zwi50dh21l8jQTbRVokj8DTT7qSfEu7DX9HoksC39cBXm7zcGeOnVbTQOF+r
lBCgFu2rTpVjb7iDp4n76A8LbMn3GmkGscBbqHDd2wOOaywmhpymLTr8SR0BRkzl
RXYKxbriptvY3lP7st9LLHN1R6tHNHVkEhS1n9Yv7ZXr6Iu33NhuYDAWkrMKq/f8
SqTsEY61hajxFDrINS6HZksA2MSUQsuP/bdyzHhFhLhNtu/AQSU8PIThtzHYXwKa
Pt6IJ5pWcDT3MIwyEIJUt7BkokG5JS6dNsW9rbTIQ5hsIKnrchq+aTQc0h9cn/+Q
uXg7VTUt/y/66t6DTNCa4BgGW2O1Taug2l+bhiIp7oCvtVbnG3ux5jeWYKwT3Z8f
odOWpou5teIpukJqZJMV42TlFLbyXPhrnMUurpRd0SwALF3HjopTLwfq3ev00KR/
yrRdw0BiWhhhPS0QSTJQoYHkUMcDUKn5uVrl+uzRnCHxHYC2ecpT+9Pm9xoMt4aK
s2p2ZXSZ61IUGDXmHlrKQlNE8A89vOscdO1/N0q3muRqXv2x0lsxs2LM/CRxc99I
IkOBBbNuIV6bxGcFLNuYxLEGCuNFwFDOfdGHpBHWwK0SX5UgUZ2qAFFH8hD85w8i
ooMMT/qnn72t3dSiuwDl0R+RO4faq8PzYldQ86PpibCya/a+JLgQ2WJZmaXwQVbw
ce1CdGttdLabrbZXO7lrQCKHCmEPF70FyuXlEsxoVpRbkHTkosJ4wus7VGbQJbYL
D6hCqQC3CzAvueTBrwrEPS3nNFqqchOPtZKyO6nGkad4i28ri2h/XuwbcAqbdDrM
SWaQm4frytcVsEK10npG9GuBwkRgDneUL2LgUxdAcSyGLF0xCa4aR/RottCnp68V
pmfYDgCpwk2LFu+G5mTwIFdA5mym7sQtbCg9ejqSu6KGXQhAvcggCr/E6xxfDSW9
UonNVrK+gj7RIk+qpIWSo9Nbo+X56ERQS1xPLzMO6yyHHqosJNRPNKX7ZU/6kwHM
Pc+bA79XB8yE8UqSGvNP+fZwM6IIdjnWMyNJg4++zYuYFfgOvhrMnvipv2UyCoWE
HuvSlLaIimx+JVZ9bn+G/3rLTKX+1hp7hY5KYASEVMAxmTteX9PwjpSp4DzYaltf
rG9dWc2d3xGXl2AeteYoNxiQzttJh2PXS5vA8Iue6hZc/6+lx2smvkIAsgIOxNh1
KejXOlJwyCEyymA2YEArx+rXtVafMAcMj8DYwXvkqRdEn/6pzEIMg985g6j7+TBl
OF24YYouZ73w0dZCma8tfTwjm9f59eeJ1JPWHxCEC4QO/29hjSTdbo/SBbd0BhgK
ytVnLjGOA+hM20g7ih7Go/vCkd2aC2DzAqjftytbY55BIWAdx4OckHRaP1nRcbkW
vXiPrPHUNzQgMkhkZOemyrayBaevbY04tYoxi6gp2zKCWBRK5cPR4TIiQyYuXaI+
cidO9GpNh92vMxNhRHQcTDu0CvBZ7AiIyql5zK44PsT3UJSXnhW7eduE0opo9ay4
/z30WLjmdwAA2jCKMDY0TLMz0mo3uMPCUhtrvRzGCsErHLZUJOl6yoUg1eVGCxl4
N95z9967pGPidM4HSymRAXXKo6yQw+8FYyE07gQdpqrkg+gav9eJN7WupNQSRbq9
iuYPU+3BGYqOPdw3cNni4dEqaVNeUxZfefI7dPdJVR7adXlAb/i8AKIInbTFpDi8
KKDoMTUXfi8JxII2eoscBxmTXDIUr/giZddAM8ETOSje0g11bUyRWJQhjcK4wc1u
fUAfTb88MMkFFalszH7vVH/hmDmyt7Qy09QqTe5xnxQBBCFfC4gX5ypXaNKZmuQq
f1aDlks/O0zKnepKA1N7QSKO+kfik5XhNjDGasP1sGzV5VRWsAM1fDIVZig6mt/H
oLYKbfz6pT0/xt9KdBJ9T9micvHhKlGVWHNT+aDRXJGJ/7GWi8T4S3whdqIUUGPo
G2eDrZHzroT1+Fd4m8lFSihmVMOaPNxizyHVtliM5/hrlKpJ0c/LaIm6cN8c29Tc
+BhuvHNZADVfG9gg9QnCclSlNE+YsMbwJoNjCCXYqW+bBMd7b8xGRd6dyHj7bpTf
81nepi8HolE1/zn7FI9DYXmGE1x/uIsNIgOkvD3BQYv6WG+5o6tWPauPQ27A0Ybp
gN1a+pE6ilOVDK39oQW3HQO8adjiYkxB/VErPmkd6CaqJmVFApquwwJsjSRubBa5
sWcsANKm1s/BSBJJUD4Z4qVdy++j8IPnMfI/7ETe0IQTh6NPxd5xD8CRRHTw8DmW
8d0irTwg39lWdGY0Wi4TUO0QTHGtjETdkhRYNvRBZfUFiOYjMICl65K35XZivgeF
W3E6hMPzpEk1xJuAG+0VEZdLrh0B9WWCKoL2xS3m7nWvYhbo9/BZtQsW6lKYsGIg
LMpAuFvgppuvOxUdCIkfjvvRkKjUmwr3EIaw/p+ryLsBkYml6pr0ghK5JoH19ysw
YIMo+vMgdOM1pBqaLk3zQ1pYgewFBHrw/t1O1lzBpIUAWr/R3tTB1vlpoDEDYdLh
7DitAcLhaHzuFrRcXbampPIBK2yYp1l8Osf7keOR96WTwv873B1Chz2lHVGQ6uYb
JEHrhbi/rG/v2c8h+NpcdBxNMJNAeiihDCxEEsGUJfM+gncdLpQ+CWFVVX55sfkQ
uyGrf2iOShyeyzbPmTsD9/FpI/Un6Ay3Mrs0mw1G3r2y6eEa5dNtA8qG0nQwyYPy
VLFWhU80vdMC5wzKT3NnhhbAEQzlM4jDUj7hgZK/L+8rhn2m6AZSFR9F6G2slEW9
KVDVAjN+wTouT9axQYPom/3i1dbYLpTttsNeJOWH5u7Fd3ZP+kwEcVL2z3S3yJ/F
gC0W5wXoDr5CBgDQyPCmNjII6OJvdLAOFNsSpezsVZpQIwJ2WKTD1AKBx018dayy
BY0k2W/d5Yfp6ssAKMC9HGKso2zZwF6wqza8gGkz1StR3q2jz1w1NELNIyH0Z8k6
jH5rXeWi0bFPYZK0sH3fOB80Sq3dbPqAU0/jW8RR99BlPepFrOaRZNHWDlLtVu7B
xsXTRDbEzMyh7c/pVWaxFuw3wKv40X9Ms/gLrzegYwFdF5YDU0z2WDvAsz+I1C9l
FGybtpmrk/Vuk+dOsqdin8Tbww5pWzPcLqVGpwMoFQ0w1gIf4I4H9T4mIVfFAaRW
Ie5WHG8aM+EgzSC2DBz+dkzIWXMVJQu1OgNQPdnkKeWhfSzT7xwgC8uOwXCPU1fd
bERhdL5QhwLiAZ+Ks9oJGPWtWRRO+1K2wmG3vASScdz0qj3sYXNgsCWb6pdNYhtI
PYWVJa9Qejfq7UyYrkw3qNa8Sb4HZ8JD8Rt9uzKxQKzEq3kfEIZ1ycMi03aYgn5o
F8k8Y775ppIniDiwkSd2twtsHXLelAYY9/xIJCmptPq8v0WjFR39p50EeXwIV2FR
FkeNeK8WRQiRVdK4UaeGG+XexkTga5nitsRctC6ZSqHVvqyO7hKNi5+gyw2dRVXR
+0JIUB8ohwGo1GbsGEiMjcQCjOkwGtThLf4Vy91hxxgfsdhO80wNweLq9Jlsek+v
pC6RVfzGkJx/dUBUCuY53yIM5q/ysoAndyAyrHMd89/ODqCK0JrYB1RsrWEaMV5o
dHVOGiunxprfGyX/55fZOPkpgvIgvTwDP1v+m1JgAehwTZU5Nbadw3z+OOg8vTcC
pGrcEBGCpdG0gXu2AqN25ovz2a5FhAoNwFTVi4hBdd1dEI7o7h/QuJGvA50pQOE8
99HaQcm21YlPclTj0YYH4YwROzCaf185AitWaSB+2q+GIi5MEGTfVqIlXXeou+iE
kQA8EzUZrsSduK3p++BVadadykuQjODSAgAnEYwRwoJJCrXKJRUC4QESTWv0K5RA
sMeBhoSgGRBrYdY2t5BGVhqU9TjoGWKOne7l48kMKCrJ728in+DdsCnNmPmzoKe+
3DNUwzoCX2906HJw6PoUXmhIHSFc+x+JRliZE6EAqPW/FhtjSfONtnJcEQgSfnZ0
tPb92DfvoBhHQhZMc8gmsZKvIG00WK8uNLEb179VIYRe2JT/w+v2H79mk8AQirju
Y57hDNEetHkdc0LHbPbl92bQ+s5eDal19vWabWj8fQhh1HowXaNtJYMhGxGRcuYu
Zn5deSaNIA/ngTbS0l2S/yYjws2tXOtA38/bhWpeJ0ySa6Puoy38VLDzDfYh5F9X
+tIiSdWRTUMzu+YuIYLbZIssKjzgi7ytxzlBo5gbUc4T9Dx/Dq+Ry+IVRetDohrT
9VlOAXaROMdze+Y0rhVz8tFwKDCy+UVA+DywthICZgtVcVPHUfZAZXg/vR56Ogqe
Te0HSVDMYDxb+bzsXkIThj1e6jQ6FBf97g0A+ZnpQPRN4havfiOVWYF0acbBFWDG
lplJ3MRrJv8aS2tS3Fo000VnKQA/5mQg8qwXI+yqPSGzNqsxHB5Z1ibZlBb1PTpP
ERI1mYMm+O7FHnJjpYKMRRLhofzSZESFJOsvNF4asJevMWzJdkVg3dwvj1DyD/0R
NjxWfDsLr/oX5fTOtcvQ6Si6/l6QcNu9tB/sNijr0coPiRAqHG+yfLzA8+glqJyJ
kZo/DufrY7eDEgkituxL/tGLgrN0p6rcwwbUplKtTJzQT+qGtUwHZ2kVr8VWPZ3Y
9d/IpbVXI2hcAvv14MHW2gDoCiQm8AebuNokbLowXN4w2LWfDV8gMpU/kjX3fkNW
WYa1WGpjOP3NqH6qjgs1uU0bGG0LcNr0N3rAKKvqcD13FdCIVys5GVDDP+Sm5Vgb
Y0JoxPyfqh82ZN5amcJjeG/TErHBYFj8YP7Vqax/dZG/8yl/bnvv86XZBmfCBJiZ
Hg1j7yMUqxVrU16Q+H8J+zbPrMMBlM81R2XhTIHF1qwZW89Y4lnuAkDGSHSEh8aX
awt0MJsCVMwFYOLPDOTgjtoMCPXhmjKHrQTA2VoiatZ95qYtch8L/fvvSMLbhiyV
ncK0brcY3pZprZ/tlzhYEFvwD6vuTZQ6/r39rMvt7y1bKsS6GptqIJjXykuiDGMd
po+1PwY64oKPtQ2+Yl1caDsaFosiVqN96GmnrHkkmHWlBn/cmw9iOmn+OLuz40s0
VOeG7Qj4eueuC6HZrIurV9UmRSiaFpjmc3Zh65PC4ptCl/HvmN4EXIIdsCrwnGvT
Y4ClMmrydKdFeRtdRhvyc9dUA2jnFZHGOHIQlLdGA/kuwVzmFjLvjYOUWmZD0a7J
27Sc5vr3zK6z6t1qPSM1kEH4Cd4EDVsWklqD9J2dZ732lB9pO6EdsEWTi+/qWD9I
a4uSRG7z8/3sNmyYgIoGfU4U+25GjvNDFLMPx+8Lows2X84tbqhW0O+0c6TYDOO3
x4GI6ejGaUz9J2hvGpwHQePt/BL3HTk9r1UWWcZ6HRleXeyqtPxtpq2yxFjBQX/M
9DiwduvtQspPP3ukt7CRYszdLeLbQ0Ca3FdkWEY/nclQ5vdqJeeKYlGQYKNRXYxd
x1Zsd1BFv2iB5s20NzE9+Qv7+UJ6/QBSSm9CF8JU3PaQtDjk/TeW+7vklZnrUmjB
Q9AM8ORGzfYhxzadc22V0/RrTuPDmiCVLEQezl9LoQI9ghYM4UVq4XjM0pmNtFZm
sxQoPzoqiEvzdqEALN37WNh13Yol9+AisDvY0nAhpXmlLrBap017SFW14hr7tUUb
SfMfeGzyhHwRn7UN+VCFZdbEo3H5KS0pzY8HMucII1EYg8ZXjYJODrif8U1EQ+f2
+s697DlGVb3/i3g0+fHmj8Gn8l1+fRjjypFYMgzIVo8R2ARpEbWC3wVgn7BShhJE
DEi6WkLUN9fLEtCkop+7gy3Ck86sTZc93KWb1/0THsL8ns2GHv0MYOEK7fPRZrRc
5GyCYEvBOl2Ox7hbSJTxsSZiXLNgcVzXBKPYzFsQeb8rZw1bPczMn7ZjzC2/LopN
Ryx+4sSqm7XOq4BaFUdy4DAd/9LCm3A9wGJrXMGV/mzh3/xqhO4cLIbIKGykFhnM
v3ve5D4LNlnc+dtD0sGYkH70rSfoOiJ3pwQnvDrGSmyzuEz8SbAknpxEMKI9RcxC
bZpSWUsVeSXzkDNF45mQH0PSWLTyoSfIBXZiOuqFPJ8pZYpoY9tjTa/FNKhppjmR
0PuVBQX75mf+wVk2WW4/eCHpXEdt6fLcMIdQ+ynEPOa2fBWUxbQN13YKQZBX9R3F
taETH0mupOfUqNhWDxlR8jQGoFBZzIxeLk1YY1+wK0FnkzFeEVj5kYooOjU5JYgS
ifNn+jgdH+/cBkN96P9/Io6QQHtmZ7btdbtbZtC7y+JJWUOdkYmBVFu+iaFSuOLu
aPpqK/uBGAdBTVOZQ3pSvQlqDsp1ROFdVUCTcQwEdIKZBSUIdSqJQ+W8s+Z30f8L
7VoEJCQRTpUAeHovcXa0354EzkC9k6yLztY2qVubj/+BQUcI1b6Q0v17+sMohY+a
Zu7+PPgy4qu457QLNP7wNYQ412wvgQQ4/74jW68CKnuC4zrH38gvAGoYavv9C3Oz
+NTpmU00BXK0CVzMBh7zvzEIgccgIjI5HzYhExxRY+dy8dbc+AtB3np9wTyqgPsu
hcTbKK9wc0eZyTLL3vvqIMBfN9x3sefrak4Yy+dqMEl/gBMCvsXMepu7Or3Hb4D3
sn08jTWKBWuw6CUPCJHevR2i1ZzaCp7KCAp6UibSCNgv0LMp+zhyhnO50n5c6h33
yO4OAUlsv6kKJMHkSN3rkto2nHe0OAsTSbg4YCoDHcA4VsSqLpxI7nqu3JhleXPQ
lmG8oCsoGQQLaCP+HAJZzLEi0OoHzc2NGWiyJhXlgxvunbT3jGk7xLlIVe6y+giK
7v5Yn+TxfH3YJSZ1vYlQkTXLVbM2H8a6Kd7ookW/p5DYSgBAOY1BM9c/Zsc8uPbY
n/4tB20RPPXna0JPVs5H12C5n+VLoQVIDDmS8RQAXqhXFCKMCUnGzC6FsU+kTyq3
wgcGV4lE5Aq1RUFi46jg1ccEqyXAk5qGfkpwWzbhAcTybkpj7hJBu05xq8lSbyQz
1bVtEqRVoVWKo5oROp0m8QIzSZosCWDp3ccbRiMJcByRsTbqiXz6ZIKdJ6zHDusc
BYPEoLBUkrzNY7hnIrH0rV7ctElIl7RoKl5F/SGZXGvjW7qC6vXqsqeeXG2WtkZu
c+k2v51858RCmk0jXU9fTozIMwe6b1TzYxk+1Zo/RqOiwQJqqraGrT8JPqkxziRQ
pPCwTCMTJsLHCKcFrUm6WQnFqszCR5pUM6h+5LGKieHV+4wZUJIsH3+8LGzGvNXb
t7/ls4ef0TNEQSEEEzHejoWl2xBRsdceWWT+dJoENCIEafqcy5y2Jda6NsDRMzni
cGlCdssqwzNpJQcPw+1zJKSgt4isBF3fOaLytFUfFTtTwsZj3I06SX7eRpLDNFy3
RPsgKxwt/uWFMSJ8PM9+ky13X/7OYcEZ0iSXI69vKDg/vpST9hcZ84hQRzzU2C7P
h8ITqfl3wZ9CkbGXh/KUN+PUDcfMFLgrVBUobpBUbY1uMeNbmjSBDSLzncu38bhM
YbXmEm/AviIqoI9EP2TmyZAI4NVYFV7tiv6qwsivsGpULoD1trUscC/hjz4s2gnu
PZheqS6H1AUUMwhz/vLN+khGnZxjALxc3h/DQqAfaRKJZIlP08iJZvcDIOd1bSAW
i9ok8E2tdinv4sVqve/4Zntij62TOn1Ma2wst3LAzWjvxfzQVh2DzO2t6CGVNWWi
HfK+op67nu/dU/4j7qFA/p/70LDLfUjhpEJ9x2o+083T7gy+Slri9cS8Oy56X4pg
OSbyphGEXmF6SbAkwujZ64wEjtqeQ9My9/9cOrI7lfjpqLr0XmCrTjV1/H0Bq1qJ
3RsahdkAjJYLHyR7xNnn7hT6gkTOztTQF1UjNhzGfbdScuNL2YITmdubUpYZ2bYX
ofm5RtMnjf8B7M8Go3l3M0vBYeRvOwzd4omshY/8CPt2px4/kzQQO6bzJ/uit/fx
RcSAWuXqS5rKbs8A7s15BVawQUeZX6KvU/EZDiOvRz1q0irq0aybKUfBjCGx9PsE
3icHqx412dVKyJJo7xCXcbq9teMHiGZY6JtyeUR0yB1iPfEJ4RUMuIs2k8a4sRV+
4CGEiR0/GWaIKLY2tmQH2qwRPp51MZaRum667N11W+lQ42tYGcvbqFK1i3ke7H7i
kf6eODdhIbAo9q2AD5dmkBFsBNBm3hsUneTKVUqZ1C8Jmx6gQt4ADNpRngkAX6dn
oSG45CEV9opXVUxmUTAwsnfVUCnH+63QxPeoMbTG3c/jLWqQUgnnmm3ga5K5YipP
9i4blM83GNi9gSrWzuEKg3VkK8fQ8SZ2spdM0Z9VUDWbFI9IQIaT68oF8g0k+FxD
YPy62oJC+m0rdCdtQqWTKsIUpneaoicLDcH6dAKMMDxdcM4EVtc2RekkFmPaTB8+
/Kr+z/jI3R369ydV0KE/Yz8+14hDta7QynMmz7eMPGF44SRQuTUVmht4gwtlehOR
P3Xyp4m//YdihvJLWVLVzs4frU+ZdYsm2xY3Svnzl31d4u2UAMFRXAvSiMxVJhFy
qXHWB6/3sSWScCtO58g5It6csAmN5yUG3ZW5a5/CEhkn+D2H/tQEbvGNtREL8KTN
2vxzZwMLCRPCRFM2fsAFW5UzvKzXHSe/EILPIviAkVClNws10okUEvvme/1MnwWn
q9jaw+eqoe3IttWXORv/ZQRC0HHec4o8opwslxiqPyUlbkMbjOZP7S5Vpgst9UAa
EEc37cuMoBy/siXt1dUFtpi6yrtv7RqehZ/vEwEtSB8Ci4KhbW42uhMsx0AfY18r
NTYmm+hWHElVS+4uS/IPwCBmFqJ1vGpa5EcQ9J+1txuEGXiL+unX1v64v5N2+ABd
ysvy3byX2uP+KGSKQjEBFuqf3WRsqauv8AjgxbR0LrsTjAsRN9QkdXJkryEff7Uf
1oEwA/C6IOIRFe6gtuS4pLWSZy+uNgSwjjjE2ls80w8UJtqbr4rEEes81xs9f4yO
HI8qAyzB6fysFa5dUYaRvaH1Tr9NoGOYmiybo/cHGxkozEd5Fdu7Bg+xgFhzGMAl
1v/D+2t7q8oOiQv2uWeqXd9gXvRiyH6cAS0yfgSNplSnjpU41ef1vtgbUtN8QnA4
SV6N1YJPNxjOisLDmsBKdfDHogUBAo7zFSbwZenZQtdtOSY5t1AKj88sZUgkLjnR
S6u6YLkkv2HmRQutTeIkoQiq+l2Zj1rcU8GWadC+o65DuJn44TEJC7UtwIpLqwXz
sQuQMASe5OMYn9OKda9xDRmE7GpwfMbwklO13Uh4vjc9CWmgwvrWsLJoJcNcntcY
g4ldEIPifb6Rh4YSXAXBngJzwbieRiNbjmkVvl4lgGalI1uMcEAJRznq9m7NARg9
6V7Mh2pSRBD1YFVKAsdpYWAe6DqmPrbb2n9gs5YAZ4hQmsSsJAr9n5Omx+mUJMh3
g5IJIJao7ZiuO9DFTjgmiwo6dUDtVcoef5uVHcU+/Hp6DPPNoCzTKs81CI2Nxlio
zN+E9LptVCYdsLJr0kI2vqte3Y4YyomjxG9745Wsgg+sgYREWB2IH4WFs++6o0Gf
SxrRgZINoiPlv4aWkoOTJZ0vvi3DU7HA4+YTVyIRzE5W0s93n7vlElEKAYUP6fpe
/BZGgLLdq5xWswhOx4Nt2R0PHdF74Kl1ZVxzDL1l6sGGqnPuwBIAvl7a9i4QgNz0
SeEf/SeIOkwiri8XhKw3XxcV227sewiyblHGQZ0ES/RiYwDNL/6JYqyLHVCM62Zd
8v6em/sLK9A3yIkX9evg5t3+IfMHV2mwcTUlmDj0cmhmfqzZ1e8ToH7/ZEOmdjFU
8JfSP5rpawM9CwnmnzL20XZg9dTaACIUd8mFxUjS/0qMcytCQDFhTx1EvvA9/veD
iv/ZYIeeq+wUTf/isK7C72A4V92bNoExz8+hQzVJlfUzAFSt3d55Op4tWRqMxjjT
esCGjczVivyDmyJNmEd4ApcKTwIV+EE+Z+f3DSCPv80sFq5phREBFKbxCE9oaiZO
5TNa8RwvD6KGWMqg2qsJowX6QXV0XJiXX1tT5bLtvckeciI8aDgCsFBfi9NSfd1T
X7o2X/n8wRoydHtfJzrAgiwNaU0/BAeecKaojtoXWEx+SSrw3U9KBqLZPYrxy7sb
2U5OTyI7Qov/I1E7cA56s/lkVwc5Sj/iP5+GilDwcRTRITI7S3zReuyL8K68lf4T
g1pdOyPMWcZa7tBWAITsE1ix1BCQ/rHAiEoW2IrOZMGDxNSaMH82sogqSLUGXqE+
bp6oR7o4Le2aB9/H7/dM+Mmmv1vctiHxvCkk4xkR9oauIKXAQXfzUMhBzK7hLu9e
cOMkZReaG15EXeix5Zc8GFtgAWUQ930TLZlXcmAHMuT4HhK/p9AWGvubnsZ4TN7b
W9SRb2XDyaQbrlAJVcvOK5m4/OXD55wnC+1IWCyz8/vr9GTNjoKKipWIgW/VbrI3
cgQtDnvqTMLhQdHgawNoX9vHYoobBTbNpXIPZ+lGWT8W4ln/oK0A/6Q0dSGcUZq8
YPpcBGVVRz+2ZETsnUej/XhhCJVUZ8QhzL9bINgpsStHhSPggi31XNgDLPYNumPZ
nRBUX+xpXP8vNEEqvpVPePcM3bvK5CB6PqTig8hEhjXEe5Ckovv8fuJcUREWpum+
nLjUQmL87Gb0fP2XGlpIAGhoIQYwekVFNlWvlFW0M6QuPI51uuJXk0KVBClQpfOi
uHrriGy7/CdSbRo2747he9Ix1k2g7oy7t6CuP/hyGyMdFEwsdxzjDQIs43XkuJ2d
10eAmTFAS+Hpz1a75Dea9ORKcf92Jh4+P8/6Ska9/6YiAuDAYESypBPKqPCSLc06
vbhSdKYH0/YQ6wDO8Mfw48LgYv+CdE/Uy1nqeK7KjpnFaaSK+oZwE+LTdR0AY8sf
ekYGB3NrDOGM/G7lO4mAk+78khiBLUBC/GQQ5wiKWrBod/Nr+Pg9/rppSD32I3P+
q7KgTtLaTrwLWruUhek6df+NSAoMgCL0bIl5JzVC1dEDdKDyuep93pgwNUn9ZP+O
mf7PvZecmHPbAq6KHo7GicSio6OFb8reUrMFYD4+PPQ02BioDVuXBcH43KyGIU1o
7pXhoZNOU0eXcFzGHlYfe7WB2PY/TF6+RHUT/5MF0bjoDGRbzY6dlpC456W4nVHZ
DyGwEIncOw3tsZ5iSiAYwJ/Jh/bFZ4fxTVPtDtK7HMpd9j3eGWbCxgl7Y5v8KtrW
t2k3P0yOIwivvQbSBt7wHiQExgs4jSfNgyYS9j9/KWS1iiTupB42MgDpAS4vEqHN
Vjj2iH3jLkHh38n3zjBnWPmxS2+pNfVdSobODhrrzhcWPsZo4EnLJFV/RGPirAwJ
6/MngbOudqTlM5FB+Xc8MvPjL8hGUe1l/SD9rWhkIkdkjkjK2xMaOSHQGS8cdT+U
2h7tYivV8cjAqoLkhHRy7SGapbt3v9PLTbbctahguYoqxGQJF8FEmrrv/Z8KV6m9
FyccXZ6EjjjyHNnuXG9E9VxZNX0LRjOfS+u+AtrpYUQo8aXOM3TGMoe2XwW4qNBH
avhjQnZGC2HXfILu0E83OtClu6GwR5sqR3Nk7Bvgq6inHXT2Kfb7AIKZJ8nGno+r
a15wAWH3EURuslrik6eIiuyD7chmXVR3k4X0truKhBZKJyVUkMY+dPMdiP3s+Bot
8VwAnzlTPLC/GhDLxF+83jtIiscKZjpCLmbUrISjCe7yOsD/Un69o0h1rJtphGkg
VSznQL9Jg31aiCiyLGGtdvj2sxkt7aAnsoi5xdq/QTTAdEPTm65C8tvq9XjgXZkg
B47AtHFfxHr6qQ1o5HE/Co1+uZ6jcTfWYX8KxSeO+xtjCeTiVOl2UEYWCJpVPiJN
4rcD49RhkHi0eBcFoTlfJ5LFldxjVIaG5Z0E8c+u4+pYVPD2Lpb15+empmlTvDIe
j1Dpw59Y08jUzAtg0CFBM+fGILLqLjBuvPvqP457jrF1YoU2CCFN6B1gKDJFhBQc
IilJEHsFEPIprwHrst1ZYvBrFcrC6abdD6V9PRFN5/rfRRNo73gRlVekf7gUCrKO
Npbu7yTGRKSu8LdHaCNxe92qrsjvCgTh0avKaAEypaeqi8h7xcuTz00JKyNffMA2
xg58zosUzQuN3sJwyB7EWnl4KoQmQVverPFawwAe1NelHulCMlY+FWy0weWPnCNA
PL+v7xtIAz0rOcI/MlxLhdKmK3uSZnurwFxUXygGEXWk/QZ8Vbc7nmgS+OMadULL
sCkVNTbTAC8F34BHUVa3eig4CAC+GeE85vAtD689hWBqQsPI4ryZCc0EgkCmrPVK
o8uOKyqKP06lgdR3hdd9J5oBU+XgAnR05aFt0UoGPQlZfSXdd8n/yOrRQB8jSlJX
fUHGnaT0AWWU6s11XUljnwV07uLSXHbIUWNe0pEuguYlbSxd8oPlQkl0dxJqgDgh
LZEQW/LGqHvIDZjOkiglnYld27y4SdGXe09Vr3LP0R7/B2cDViwbQDvqIBdjtY2q
RKa0kSNyzkNnzXviYcRWZR8XR6vyoYl7gDhvZYqkaDsCgV3noLE83SOGgaP9zxm/
7w/lQR6CdHu6kOamYcNXKfiMMfewdHOcyiV6brOGEKeS0B3teVuuBsy9Xqs72Lmx
u784ZdHlgRINlA70C4hUOvDQuTbxayvDakiVLs1aqueSpl/j+4Eb/nCqucOqGEV7
z3cgwkRFJQX+OFHISFtB/ydK/L+NeV1jsjgs37ee4vO0dchJ0V8QahpbGdKkGfmK
nqhh/YDcpyOqSIJAKSS96HA5WRapHWiAgmunuVYg9E/QoOSs+/iqeQj6FamfOnPQ
jZ2H+hqstyBX92nlBEh4jxQDQvaAEmorVw9cwgsd3cMLinwPf+tLvLgRA/1ZBwfd
gPTy5q44M6zqOpAOBr/QqbfETETqSY7XMks4Y4Yjq0JBBmQwvyiUXS7obfCZsC3P
froFsnvpy3kmpYIQOyv5qZqi9uyAtgy0xXbWHuT+v4x5haum+7BxrELwi+PP7B3s
7fCNEGv58KjNKaqUVQ6Xn/DBngd8Rq/IQqGqqztjj0Zjo5UzhBzQ53XsqF7knQ6C
qDraaRB05w3RfdjUJXRwO2RtxRtczCH97rChUq/b+j7zPNKhjj6Yb8TRquoRsLfk
TKX1dnQ8YJCBsfXgW7GlarUpAXY0Yk3u9fUsfGC/7mO3yWsLT16ZnCzU0WfCS4vl
eehUAuhWQ2jYUA2p5Iw3AZlm9gh1HwJA5fDw99ZSgCD+bkXMPOcTEBDj3v7N1RVE
PrkFzonC2saMjFxkrzLGBIbaQ/tb8dEyFw9UFZfCFAdisizPaEi3mggWSKfrp/mI
qQmNK/adlHI82K1H2fkg6wxEffWVj98X0U2iC51HYccfOYkarE85lv8optBvGYiz
bdKKmg/97FYgSUi9iBnU/IiXU8AQfe6P75naAeqtHT84D4b5g+3UBP+m2XhBAwr7
iylsIgKDqjZT0AxULX8SveME5gDxUW3gbLmvPWs6ZC6Aj/2W/mQKh6NYa0iR8s3C
KxN8a19CZdwg6j9C4JmCioR9ornpbP/K60ZKQa+5dTC4LH8s5wryMz+Hle6HzJID
XM6z10+bx+kja4mF3CZGnK7tIWobcDjHhuEu6H0ylHHN6ef5l9eTrBA6+ogqsMhl
ojoZhWTbYXxF1PHYFSIvJ5eKgTabEZDqeBBxi8r0Qt2fTuswF2iTDogoxSr7fzDZ
uH4+u9iPLuNTC36Xzd4kRvnnlXMWLt5FiLuCRHhuu5FsycvXV792DWjjJ8AJcvOh
NHYY6ppqJ0NZaqYvhjW2sS3DVQ5AeAIBo95dhNQNxXMp68tq0VRdfOiHZKr8HTVh
ifiWbOoTl4cEQVMoNaK3R83e8zIN3eENyyUBJf4M/DUxVjEoIOZnDW84ABkESLud
pucB+KQVsyTPICfQvJ45DFX5Zysz8AyaQ7d/gzldk2AtG+8sCHGyowyQeyzXR2cI
ByRataxNdalQHjk+xRxG6pia/SByRzUkyTZlcIh3JlZKTKKCvsU9mY2uxM33OkOQ
o5scGhdeoeWoIf5Dbi08NtV8JFtT959llhXaMYGNk6oOJQVcXBRHuHa24024gM/R
kRl2xu0HAM3fe10PoGs927aKsiHJwt8tQD5Hattpuc8jMTklG5M9GdeYYUZb0376
8STDMCVhOV5xBiRPbYe3LFPIVHZjl2YAPagV8DB78Vw4yfmbEbo8c0WQ1McKFFZ6
KGhQW5PdTQngzqtRsioG+Ya2tJrm0DbS087QwdwsJlDpVnh+AnRC05YoBSeceOUd
XI//yGnDunTBDU91BvD3bAP431UMvS8DKFbU6nfocc6buFpAAcIqoE61kLerzfiO
qdKmqOGvYzft9EdD+uM1W2T134tdEuYkZFoz+TOJiIA51BGC4NCjht32apD23O3u
m/hrvK77Jet0231y4UuqGIKj0L4Qrzvr02/X8pURr0WLx2aHO7gkv0hURFc7A7hK
sNLo8S6xKQYmFXu4/u3HP1C6k/wmJbwpp/Zb4zM2hKma6Ro93id6LN5bUtmW/ZJL
UoYGdNiyj3AOtV2LsEBK3CmTAidbqGeOML/VuOLG/iSq2BKD40kqDzR7N9RvZwGX
ep9cqmx/rMRM8Mj24LgVu+XLAHzw1tG8R3BmttVJxtgxs/BlOt7Y7XPb8b4hWHyR
0jG/d6EA28P+Dw+Pd0rhVVnZSfQ+5lCi7qyFE0J5El2ZaYzCfyQtCogAiDNTyJ9Y
UChiJy/06CVrSwjBQzX1ML9ulDBOGVUM+jz6yKmJQ+dOixVpnZ8b2AKxv0AVH2oV
hFGsFOJo9NxIXxuEVTHqc8m2QXyfN3DdBgCqVyZgo0TwEF/+71SVmWy858inoQW1
5CUY+gqqiWISs8xr5T2dZhbhAUzM4sz6GxZNvdRyPrKFGjUNu2TNl9JHXMfscwTi
xHqhkqKSbEQgPf7grumLIgPye9DLc8p8x7t10YpaRyQsy6AcdWJCgHe97ZJvOgzj
giI0vqGQykvlh3Aq7fqNCOYk9VMXpFeMsqZAgY+M5pDNK04RKDqn57wTvvH6zFLq
UBHHUxNArFXL5jXxpOjE0Br4iI1nqMUKtuBZbFZLMiH4pmH/RYl5Cluef9g9lmVf
OAC4/3ktDMVUTIWn7MU8ssGfCWvp1ucXPO+WfWUHVMkYm2v6LdOGkUN0qVJCoRej
gr/9nQNuTmMvQT4E8coO2iEaWdX89VmrmId1W19GJcQYkcWOsWNbU5WczAOfq+2A
MXo5QjB/307m9rs7Ohpox1YdCqKMyx9C6vF9DADYitpscrwj3iU+wKSFnbHenAgU
cDDrav/B7itEN8PReyT1p2Qtw4MCi5PwNvIXUysXt6Z097uTGm63u9+Kf6hBMSpF
YmXSm0PqyOTnbUKdWD4VZKkrnkSvnHmewMNtssZC4yxiCh2rxhaXBpE4prGsFPcD
cL0KMnS3wS50Ypdw+PeWNAPsLBeThC9C9jWG7xp11tqYPSpx9xeRfhPgx4WySrjG
oL8kXjNWRJizn/n0rSC67q9EVJfbRpAJbsbgeAM1PPuROgWyy9JsJuAiPAg7lVOH
0veOwIxCto/XmfAuP3EsNLJ5EReXNl4qYC0QC8gsqjaXGBTRN72x86RQ45zVxU1L
rZhcEJ3ypImT5P6O6ML8/htIxlCZa6twNyqv7//t0XL9ZnIl50rrZAkYMUmK/p2O
VTa3r8kDod9omhvYp/KpYJCmdH+roVxfg9cfdh2J7Kq1Yqq45i8ghVb1W4nRtwz0
E9wJ6bVRfCl5uUw4r/a5UDGG5ub+PImUk/f2SMRsyYv1n7ajfytRMR4gixsTpCzM
rU0lYkekThscZljB1macL87f2Ct+12H4yKo8CERMHVZDWCk4C8Q9ZktdVO7moBai
3wc2WpdR4bbfzSmDGqnXUxCS1AtZ4S2SNk8AJoZJwnbJjLheSg63sPVV5uox+zOo
ToX0neELl0f+nOhgV7ZbYXlHrdecLbM1A+dWI/T2tXNYmiHbZVoGJdlmc+2KQAFC
qOv+1euzztI+aYFgpR+fAqgtuul9cfKc2m5wbMelR9PEc95wva5XKxGPArMEh9+Y
Q3YThZnzYkwzh21K67r2VWx7I99Ovu36JGfFViDEwW3d/8Tc075TYi7kFFMyGD0p
ZmvOlHuN5+uLnKDLxW24L8Lj47aPdgrGSOYG2BHLenf/fsPV7r2F8RljT3r+8f9l
PaIFQyMrjsu6lSaRlVUl7Hne3EOEaj9O9GgvIKU+T00XrK8HGnfHcQbTNy9ovnr6
GX4pEVcNIlAQjTqkEHIYEQABEdbLFv31RnK3BuNzBo13MIZ2afmX/LqGMUMpKyuW
hmaZTfuN21wCk5iC3Xd3xe60HL3o20lkV9ZD9Ysp6mfWhReBv6rvSUUx3kCsF/iX
Orabne48XdLIBGxXbzy5V1EwOLzJsUVyEQRRmmKWsI8mMjRxCsrwMbe/uByIXVI0
+9cOrr50XJVoeVQrjP0wS2xvccezOOXB8w8tm6pmOuoHtEKSbuDAZe2Xf1C8nnyB
ovn2H1KsyYUQBddgQwlxI2/bQa6k4DDDmaKEHRXhM007riCHrzfr2ZdGofl25A4l
cH5fFcoAcgztXbBzF3N4KiTM3atl6kofapTftWEMGnys+kmDi84MGg2PoNf3oX2m
157jGfKb2MpR02eaAGGBIoISiu4qmuP1KjAv/eK0sORU0GU3ge0XqoCYyqBOUldb
z9RAl3cJ0lJRGbP3VhdfM7VdOl7/iDPUCNUZCBfxjHXM2/9IzdEADMvZQ1C7uW1R
TYFRPe9ZwRKGS219CIpI2BDHJHTMcbcJ3LixwPxc+fsop0rKhRLwE/1uOPURrgzp
Sjj3wUSt05JQiBSNbxCDjLWcD6GKH5LN2kKVgTeVojXYxyu7Ed81QnU1ezcVPYIX
XUMFsKENZYf+zCOoOj1IzmPiBwunk8tP1aGcRjL3fgqw2aB9tkLkSFr4mfq3FQoR
KFl67lsadu7JClK9iSgiVFSGC/vymb2gnh2xmOBo5XEuISsRrMSPU9+e/+WEkldL
JU3AuSse+mGukGtbL0TuT89RUcaaQiljqxQl2RCzy/WtziV2CQROqJufoLT0ff2Y
9D/fTbPQ7ND2AOtLYOPTy29Vo4TieNycYnV0Mq6u6GDHuPXOOCUg7eRA3lkZb+ws
o5U3gXCjHajceif5g+ZFW7ubon2EkOqBOfMJxV0jhJ9lQDfhWxqTqSKx1pWylPk5
8fh09NNHjy6YiEH564yforTwXuk6jxkfGYtFCBJ+xm/NPfFFGbkhxtclZlX/vg4B
ArECDjCYXasqrqYOUc88dvQdneAXYjro0akzXZT3UsYg6faLm1FUYl1af6yE8KHa
o0TTvj0gxde6m6sCxqlufdIN6RK44zK6HRRqDaf5oFpvNKraKbPuLPDhVnZzeIuF
MBqU6mhUT9FCP4gFTkKgI0l/GRQNCR1x6UEmH/Ocu4wUn9NhwnB632SlXk70nfkc
8M39be4aqCksUdgBSKq+SPZWZOfAuIn9GrjUhYdNtFXAS6aaJq8oAaotMzKOQ80C
ZqCfv2FiyhT7Q7nPyZfld6AXnBx4rNlPA9mcG5nLxfN414Q62tSr3bMAJMAW71Pd
cuwykAxngTmsvviJkJ1AV6LvCU5v6JZ7xW0Mmhy46HH2vAlXf+/Mr2ckxw+usz7D
J+8v3wIuUBOAgzh905XTYhOxGC1afToLOTm1PIMBWWrDh9ZjrZsc5YbfQu71uYIR
76r9v4rmG5jIY+f6g87rjhmXsmHViKNhBTXVw25jZ0orBkXIP0XWnp47ITGhC45E
9OZwfpnR7K+eDX8t2xBGwOp6JuOil0Dly5WA1nve8KAElRt22nG72XkDb/TSw+Rn
oKm7mwvxiCttYgSTsk2S3Z+rlIKrUtbUJlOT4pHh5czVPMi4NOzbssL4MGbKEhjJ
Qz+3NhHCGms8cpKwkth8c6HLVp8B9dN076AYcINmOd0coHMnDBbPtFzw6QQw2UUV
Dgsx3rHTNCdeCyXDEVVYn0t2fxh1EPeYnRaf3Y0hGB1O+0XABwqG5iZ4b7M2/upl
bvobSulxCaVKzlkRMzV9eEeDx3y5lfBdpnlOdi69FBV3WvwNnr7/0lDtFqjreZUv
NwxN0UycyxnkfPap5urzaJyB6tmBWZsQeXtq0Xro103XB/vtaVpdEVISPUTLA32e
uo6oP559aj5bJgjeBLNxSUtUdVXV6WEs0IC4/cdcRVrBF8COjbdLI0kuybB0QQ7I
BJVNg7YPBlCOlmx4SoZB+zmfmmtLo+wuLVtn7PZxEfmcUZrqQvJNpXjvbM9IFwXn
Ks6sVnPowDzQQjwzQKUdRhuAWqn1Gb5DC7wG6lVMJpub2GWsbZkgYQReRyt+wYK3
feUMryxYTVwjQ9e9JsApvlTEVnYcOGZNKiNEU0VvSGQdjwcJdlpCqAtME8jCRYxQ
7N4c9vOoZAVH9q2QyU/etlghlTr+pMmuIXzmn3tda7nsYwKrTbGFtbhTmz75PlD8
6zS/3svmFDHIEw+jja/Ix8pylhFXhzjYZqaL4xh2U9XJz30QWoWNPYN8l6veP9aQ
Qm6Grs59+KMXWS3mYA9+v/PlKMnO/XNnihmkW/2UscuY8joIBzvLEq+wsQ2UMs0N
0wqR5uf3ZFRKkxo+K0ZCMwVDnmOgAflcKMYsl13dMZku7WfVx7XbCW0gj5UCLAB0
YSdfu5EwG19qfFdgEM4WjZf4ovajvYPy/Ze6gcOrqCCDbfz3JsKg2XSSliUqCkhD
IJxzcqct9af06T6ghHZfpZs/6zdeahPjHcMscKRV97wUG7yzC8KNuxZ277KB7o6Z
ekSkvl3h8rcuG+hCI+QZGl9C3CYjMJxo0mtcds8xSXY3ZHxC1Dju2LR1AIMt9N/Z
4IaPWJrVYuleTg/1OVEhd+EMLYH82TEXmGTQBJuwZjOmpxWZnbrnVcouiZ9ievHI
w9qW7z3v5HI9s6H2Nwkh59Gab9IWAcC2dRfVKVbmyyTbjXQWrRM6D4hB1uLpf3cw
A427XKIasON1+85IiAUQLT142AWTGHNEtaALffM+WMWjiRqVN/Au8o/wPM/tsntV
41ZXLHrzM2oVVx3O4yDVyz9ia6b1xIDGepWLQRbyV626JN/p2DXbZbzrNjpw2lCU
fGm7jUWCTBrsOU1Lv1hEGC4g2tzSLaMmbZ+W2e+X+ralJNSjUnW+YKiWTspiv3IF
2HZ7+CrpDS6rflvVIXyHempSowt9TIiSQMJN5egXe4ZWWPdFy9R5TcDNhiiXOX3w
+BihsP6c5gGxwZ5xxjcZOlh9CsbH4QyV4pt8KINcIipuRZSKbckfKUiXqKcmawMB
wQFAD9/PzqWAh+lqK6F2KCg+e/Bs0ZEo6HYyrOroepUc317An0T1de61SIZNWnZW
ryYZ5rgWHEflv4w4LadSHyjsI/JF0GYnUJ+XtSpcON+fTMH8wo8XQzD3uEYXOm26
Is/dVXAiJRhKw+rKsPKjBaZs09d7ipPtGPru99vRrBYsYMq69ilbXpN4ZuhtQ4y8
VJoD/rY2ci/wvdGE+szqNYHr+ZmK2FF5/LIOB+ViKdWvxkk1dgmbAmzxL6wsjQ/R
jzjeJ0vOO49KOGO0pvX6NZjSGwostoehtqHzkn2SQbshIWU30Nl7U2ZiHl9xVwxe
i744aL+DEHJw1r7qmtPcuiSB6GSW2LCucw9YuFuQw6JLXxsz/Au49s7kZSxjLahe
3fkgGf326xtyQG3E17raGouV6O9Hzbljno1zpKQ/0hvHTOgeEFgkMkVuge0uZs5V
m9avW9ZFpU51hnRivalRkHWx/W2rzr/GqyjshY9fwi3U3yjT0E0TkDOz5/1QTdJj
ujVQ7N7S/zUATyVB43u1qtlFLgnGqmXeDobHbil7WTC3Y3gkvGqzwBJ6NIKHaw9h
wSbbZiVtS8y0hHkdFLAfAMeQ747+rCYxYzyjOHimPKo7EJADRVQFWtlE/s1IKFxq
2y6Z9m0zcHOPh5yX9QN64FuZDs/5oAVlXi2Ru4M9DjEFn6F8e+FzQZq/eSMAg2sd
c2y3jAOvQCDCBA6KLJMbxXwL59fV4uAj1yCjfx8Zgu4VANtR3dro8R8sUXUV7dYh
eSofuqyWPssy6hACkAqxHrFKPedzG7qCS7s97tGL/qvywlZhItyXryakm+XBE6l5
PElGb5oIW1eqQVNcx+I036YMKcDp9K/jXEu9bzjhJ9i5/D4t2rnlqXrsiI8QT8eo
j051dk4F9MaztV5X0vHgqD6bC2q9KSV5ozbr637JU6T7rULFvMhhdhIjmZslUqyC
aIz5XsomI91UKQQlQl/K1iNpn/yaDqecPQIcdsi9Chp2A8SEhB4TCXWtoD/be2nF
Mo0KDUCiBUVunc6r5lmfx2Xa63sDkbyd3Kj3gPtrgMpx06onRyvkRPdvS23htZHc
mhaj3+TPgAz+xEfdv8gOAyFSiJB2dSFoAnLumbIeT3dCO+zVC5yWKQeGcHKUBd2q
GrymU7h1yQmng6D+Uxb+nH5TEBDXMVrytwkQNPj+4RekV2ZcyZzxM7Lv4rpiC9x5
s9/3Kev0OKX7Y6XS7nwW3U+5kRpwHRaR1l6inCJwdEsVFq4k+W3siGkHz8C1qeH7
O759v9a3U+eeKK6EfCwb4+ql4yZkbSZgAfEjaN83N5VjAbeEsVQxcafVE+iJ003x
FaCtlt1NGrenezUgdFjw3aF4EAQ1PwR50ZlizfMTc9IkxrjDByXyRZZwluAL8eoi
gqly8sQuWv5c+cryxnNqx7pUUkvxPWheYw4Rg6yXckcK2+r1wtxuX8ECGRtHh5Gh
cUiGReaWGXyb+09eiDoFwMf03dh0W/nA/Svd+D9wvid2zwgNa2+BrSf+UbKQlKl1
SbrA7ZGuGzDXK/uHd4MWnFRsWmldQ+xP8k/5lNYfeJ09Ky9VSi9r5eAVXshP/Dd+
eRoLyXhixSy1o3DRN2ZGc6bnEudDRQqFJdx/qq+PdGvmRrluj8N7VoRKMSn91yyy
WQ+REK7Msta+ahM6KF16Y7vkIeD7Jn+AaqdMg9bDFIIf8XAy7ewUiotN11lwFw6B
9eRr5BAOdyTk+1yeY6nqjS78GuHInZJIqKoYDpz9A+qTwjDLfQykyN9k4JSsBxHU
SQrUUi8fVdvdczmw684g8EX2Rp2e955UHXZb/WrI7tJqSm5vFPY7sKhK+HUVUyiY
x3nUT0o312hr2Ttk0S8RVeUaUvtclLXNFVS89yUgtC4Kid6dpFo/UmI0M9deuBzy
Xyn2Niz0gyFXwhozjHzA1yt3IEbS0cx9wK8Lbq7JOdXjnMkwZSHmFOWjsnc9DdsZ
O1RQmHNZ7k0mF6WK/7Gso317QMelbLazubbqIIpC7iw4lWUkZwR5vpRGw4Yhy4K0
mQB8wNpBxqxq9WtridgLITHqHF/YL/88CgZpewlK9rSLHq82XEKAuAM272c0yUjz
qd0waIkeSE/b5RBJoFWFrK0dGZpiyy6B0gOeNDLDeo/CaU/2xzOIqFa0ujmgjAsh
EGGSemfU+iQKCs90h/CNiHHY/9E91nEVOh97l636OED40jJ66bjK6oAoBHTGI8gt
sPAbrjy9gXBPVK6ncaSIiv63X9DT04gm8wA1HKhRhxtlVlKI7V9bNY+SzwgwpkUn
SJK4EWLIvFzeXi5JYjj7b3qMKSKBdXzKwVjMD5j11NzsAskYTRdGIZpb+dqvXdX2
sEgSIbTbcP7iUKw6eRjTpMU/UnLuX2a3LISRI79FK/0IF0xpWZ5h30LinMuBXuTb
8IgmG7X0yJThInEXGurvxETyfabJW9lGrE0ueYChLFi5bF8M/cM4ufGuOu5QvF8W
89mRbBDVzy5S69ErS5N74N+zOLoye+tjTTv4uTUJ3gAnSvPq1y8LtSNmAykUFV1I
/8r7iANpqVhNTPWlAlz1uIDnSjkaMA7USbhf3nR7ugzNGlQ9XhBglKJ2FCkuk5D1
0y/PQQ6TNysbyYH47e4NPQUh6AYoNfh8/EDTLff8HlKJwc0DQOHIRroSHDWqxy8Y
F2DIP0wnlUWXaArwXi3VISE5I/9nQqMrgzphyhkcapWvsX4wUU7bJicYT0AFvUn3
+wzYB5q6rIpH6slHcd59ixNsD552C1M0kt+8Hn5lsbJcIIeXI3Jqdr0vhsNe9pjQ
+OuGotZjObvCPX5TOJP8/VI8Uo26iV5FZjIzg6nBv81xjUC2yU5UEfVkRimI8hH3
floR1uHds5oyvFNnUYZNcIMPAf1AvovYKLYTEOLLbaJAe1fdqze10ILu19s8UOSU
dA3XdTLl7cKuCdNkoCj5rQGra3HPtqOLc1w5qep5QrCUqPYZZzRkAE+GnbBDqAoI
ImoQ8qe3MwQE44OtmzLqKQxaRoZx/NSkH947MmLASjpZzv9P+IkN2X8Kw9cRESMC
izEc3y12VF8q/os/1Re8Su4q5mR/Q7YMcI2N65fY0w8KZI2d6mlnmPNeEd8HWtTF
XaCymRuw40p3pLWRXx/TcN/N4sBlIm/0vnf899mjMtLW6jqjOS8F+mZ837kID5sf
gz7Pv7tL3f3dwXG8oD2SiFRTig3Q6ryqucReiHxMNz8pkSRxqLchk9coNxCOeDtE
k26zq0dkTiibQa/my4dEZZYqUkHkDPOgqb+uEaUokPvau3qkogvZFdU5Hs74fwof
5lGJMFRr9zgLsT94ArM6YkEIx6QsD34DUR2cm4hfvOUm4xT2iZ+ADCQv+RG9UjeV
eOW9w6Yu27po0rwJpyCd+lf50OtVrjFA+yMhjhM2Qfd8ao/cE7Jw6GL2h1iHelcT
KwmVLIKqIY/PxM+KeydRLEieI07zhB8i0ORqRJ+uAbHMtPrw7w/ICszJne1UDyA1
Cd43T12jWTFlOlHYAqXdCU8s0vsUwwMnCSAyWXYDL15EoYNRbi4eFxQJkPDy9BxU
8mJlaRmefL208+dP0G4FnXt7sr3gAArC4iM2vLxGyY/VA9+bIGO79K25aLtVxkCs
sV234/JfpAxV6p49GBE0mONYCyCMw47imTBvFg99yQFO0FsIF/Y9s0VisxavgvFX
cPkqIJB+J9X1FYSMhzTGj4MgQOTszITl2bB2qY/UWbPj9LLS7nl1j8O2KdbALIfi
R3TDPh+zeCb+lpHsup+r1vW1b7xLYRZhRX4izgsrherNoKdeXBGRz+Q/9FPQqcmW
An9a2K+kQi31bTEuIwzCXH5UhuEoiUx4z3PgPM/HKGxfbWyeteqRfm6RXK9rAJ7D
P5y9/ZOaGWTttwLUsvI0KFwzfi2CaoprAE+NmXBjs6yI8eRGI59Yw5Chu5YcrfVO
z0I7mIqt+8Qy9iNALGzPSx5UxBPI2UkBafa6NvPfY+1uO5H25yOFSWqX8dHY2Y1E
xLNtduWo7PgCen25orcFFZK2eH/q8I9KpmK6JPouJu8Gu5Asr5QeCyiBq7lN3DlW
QO35PQk/EZ2c6aLS/perJCovPM20F/L2Zn1ueNq/QqaIGln3bupjE9mzW0NF4W9V
zzVdQK89HYxDy+IALycDBOfFmjlGzO3Md5sQt/G0RLSJUPz0AasfeyBxAb/LsH1N
eO6Ur7XXMNgUjH9W6jfKKrQNSW1zGpMnmKfzCrYzBqsLQDEjG2U+8P5rZwbfMsiH
6oLoiD5WOSU3XZFe5Cvjx++AbHi0L7UdVAf32BuJoZUmUsvwxumK38qUmyeGh3+w
UAh1Lex0Y8cRcFzC/6z2CkimfmmgEy/VhPw9kaTy6+AZNWtssm95usP9QJEenkPa
j2oiD3QyGyOqYQt7L8k60JIJPvVZ28fUuUtUjkQj0nnY2gHHWojqfhWBdDhuTPit
OFnh6tNxPvIIaucaqwi1rXhf4dlPc4rtWgJwZLrhqdpuYYNFv2h/9pIaxpa+lYfO
I4jLPEZwb98/n05H4vMZ7dk1qgkjxTFAc4895bkrwdxMjdDFiE5sVj2joGxmYq9B
5yTau3b5TBpk1h9PCp64TiGtXQGPjhkgivWN/SLryV1hXM9ObLMZTWhwpqtmN9/D
nARGyOEPEi4C4liWWYcOOMH/N8WIOxBc+NsSOEMpuwKIQkzLwvsL1niMlb+3i66x
DsY9OwZFI1p3iGYT1dy/tL0rj5uy1mJ7BN4vJhbNTgT8mSN3W6E58bVl3riHzuox
27l7P8XmkLqr3XhhtPDGPnj6bMznrP8hiOB6RT7sdaCOP3pLwFow0LboAhPxRl04
aPVHCtsfTl3kBBuKHPCD+TkUx7ni6XMUOJvdf1cpE3yQRZmBorvltAzDIF4IMGra
M0GD/SiDpdqP59eEMX0o8GyU/aezDqut5nOlcAt1ynJEGT5pnQJs8Vmr4dAj4NcR
52GMGkAcBmTyhTEONRFZ5OLUSkow5p8imb9knk5vgigJapAJgo8EndjjUrYH4IhJ
Tw5PUIHHcNqvHXmItchwNVB60IsvVtcZbfCLUy1nyUPtpm9MpSyJhlV1ccO9bYZt
0KVYUWS8r2mAFGrknKCYniHGm7njS7yPbGqahINhqXTxKhMfzKFu+HmDV88iqtao
abCJ345PVw7LQH4+dv8XcOaule2Tr/VoV9EtVj/Ykx3xc2jhf9OVcMrfGCCrVk66
MiLhQeeBLUwrlvWMAkkZ5doNR7itKsxAn4AymUCVVlX0difpTmCQHXgjJrHZ9z4z
IUHflVNnnF1ZFPLcgO5apGR+EpdXVVQFBcCLAwCJO6kJ7uf5bzy8AbIGMJ9qslSY
p/t4tbzTEEXA8dnxrosaIne9A14597bljAp7E+6amGRrSYJHqm0baH1iH8iUqdyp
2jslb4nHomeyLZn/Kt1MtBwsKrfEtJU7ZUykiilXEh7rn8BrMTg92oR7co920XOT
rGyVgXInmH49i0Fl5C+rOpWO9rZiiuXx4w/IaefYNFuMJRaxct/Voda+5jj7+5Qd
TVQSbItwsKC/qFtT4fk3+GOC7BYIL2y/s14MhdgBpxTKFaGt4VWzMSxyBRn6bjXc
r7qMX5MPHfraMlq4L4KZl/24J2S6EkjnNjXJp60Ad9i6IFgQW+Hy8sgO8rLeWADD
eMif1utWi/XSNwUFxI+xJJXP95+6OpzUoNsEfnC9LLz6LJhR3s5UMNKQKjaqwt5t
rQzZFuP9Q+iuu5zYSUzI442xSmmLUdIDv7ss3mp4L65XZswT1SgDlPuOnwCshiY4
uM8kBYXYBvotRdY739aXIub0vVBEMYBcEQVW21Cfj3HxsnvmhlAjHY9La6C9iU4D
YJjeXAsQv5z6T11R3/fuMTqT0rb/BBUvu5Dmef2HA0K1yCOD5549p3PVQD+PTs5t
scdG4dGLo+61rqHeEoezE9zsELbET4349gZzr9syi1+SdKrGoyREepnWBKCUthbi
erN2CAUaQTVCnsIq5M8gVDJqIQNsM3YexopWDg4U10V3hz+MVXejm1KQdNYzBqbc
FdklocJdPfTexJE5g+50tszxVGuLgOnRY7vor3TCwCn+SPrW78GIyUc3Qkw2+MU9
k/18sC3TjA6YgAzFNy43Jue7pppSekg7X2xIj5Cu3XhziDpDPfM7EKJGg2frPY9N
eazyo/264fJFkjG5wwpd4Ew9+3MKbZsQXgLYYDoeealoAYUY60PAL/jQtl3Ums6F
vwuFMlPb2hwcwSKWLVJy/Xu+msuaA5p4+i9662oUNo0W2ynaYSV4xt6mn2TM7kfX
rmJk9OIPZSG9ArlZ70EsLeue8M65m26x/WiZ/d3BD6SrYlfCHdEpTTvpqXWZ9MCa
dhzisv8U/TPDhtN1tNvqL0qd7LmdH2r/5oQkHPnKrfp0ryf9zYp2Pwa+wOYTwvmJ
0ik9DxVNm0EBI7ON6SIRS082CnbUlkWIQWnVZeU9MtT/1ZyWqn2j6YIrnZyk8whz
BrGgolWEE3Yz2bVHEiEpHaEZz6hB7zbLcNhGgIWHdDVwijsyiEtXWzmoNEoXbG9p
4YT+L0fMJfc6zgi8/v353RBJk+LA6Jv2xddaSZ8bdVwRz+JjH+rYqFQXZp31JbHF
753Hpo4loj0IKcScsIDE+sJmQYUsgRsmB0wuFYwe0EjZNAlUKExIL7/gy6Zob/Dj
RAOIqh+nP65JKA0S2YoFeG6WEayIxMmt6svNAG9yLYYXmz1HocPpZDWt8qjWg4BK
XFJJ4m51n+SqkaS8tkO+k1eCu2fmPvYlvhRfmarutxzzPV9DRY04VeATEoirF+sZ
grFZsAWKsOHexgd8z9eFcCw1bxH1YpQrBhPVsaZGTczSDEUx7YBCagsWYwrMjO+j
qz7vfXYCf456J3qZdS/b5gwgJeKJZvzx/RhUpskaPFbEWYpzsnUKu9B3nhC6vzLQ
CQ/g8URhfCWhxbwpCM00i095AXdLxZhR1t1nzmkQvBN0oO8rrIVyGmUQGCGALWS9
2Gr1NF2KqNaORP5go8/qfM3D2Z1e2dC3YaeUU2bbpJwn5kf15t5bn3567XZcn7ga
qzUSJvf+iHYx+J4O/OJOw53u92XOfFc3eoqqUVWo6Ew7EdR0IVDMgqibLpHmxxWn
HX2s2fq4sqOZiIJ+A4eS9UDuw2jenH9hjIHXsC8R0L0Qq36z8w4u/UK/pWYoTeKt
h17/A6jhon/SixOpghVTGTpFBw+oyKPnp7cd59tlRjdSEJQa+iZupSrhj78qdpZk
x9Y5KowQj6r3N90kficSmlPBTdCVAA1M2C4TgVSGdJXL3cBVM8KoVwAU3rQ7KJSr
9/Zrl7/X4UfXP6i9wAlSzv5+UVGuoBRNd8yY5mkaJ6Ro9c8WaECAhBprUjjuyO8u
KE01rcA16JJ1sxH0HjkcdFfZzrCM35Y988M71rMNBiiu+Kw7+cxbDgXv+fadfXm+
8ThzskucSc1RCgUXZ68dw4QssfiztRQ+Q+t3zmDtqx1XiXln9DuJLe+aP9hypBtJ
hR0X0FUCD5S5/MfHYT3Haz9+lihwhm7f2tjCFVOHbepz4TuV5yO0Am/ZzWrRHHSk
x3YXoRKTCSUDw1SQj6214FYyAPT1Cx7DAqUqzvcrWjI23FZlDPG81Bw8AihCj8kq
6oJ7R+rdG1HdxG3pa0d2gYTb4+S/kxkZmFkQHX6B3WXxSubJC/G0FAhdtHWiTC5m
wylVcLvajXs0gwfF+Oe6IMarAJ1BWyTgZzldb16zPSztqtbvLWpUCkQdH5va+lMW
Z44o3t8Ub5gFCF/P+0KIbYhFIUHTyS/oTOKVfbE6r92tw/4Nzs4BozeLrSIHMbYo
rl/n2PtkqrQBmPlhjSTvgFUxte/BZiIWXTr6bKcEVq6zo//jjxfqZk4fgIOlwPd+
ODS2Dz3QtstMusUgbG+K1Dp5lbNZ+3Ko7HP+kqosn8EsVm4o6FG2hsSvHqtaMCP2
M+SvSvg1M0+MSIyn+P/znxEuoBuxz2Qs+5SrvPeNawlq6ebOBgxtUKbFnzD9ot/R
78U3y47TyffvIBxqPB71qOSQFobJccth2p67KuLigVAfs6Zcf9qdXwb3hIkmeojN
jcQkBBwmXwQyIKWSFqrQKMQV6sVWdvVbtHW2lsm+UeWOHbyzJlBb2OpTLdEzZMMC
FnNfAD0nCCl24gIeU4NJwX9ZyZiIJmY32meL9ttC9ApG95iBtNhIGLGNvSCbcqjB
A86sS075e67H82frQypZwve3LieS6e9fjG0fuAoENocoC1Ygo3KiiSTI7KpFdoxh
Fv+X1iIynEg71osWEgi35Fm0yp9foDWNUQJI9kq65rzf/Qskw25GOJxVZtSaNbbE
WJcnW4woD8p5aXhwmSJm4KaeS5oQ+Y4vXZJ3EeL334/Bh8KF6ywtcp2YRlp0m5aA
ZmcTQvxdpDMwh595g0MOT1pcJAkc3U+u3uyx9g4vRwvHmUQX3deHFljRApAtW66L
6rnM+53tZnn0WZDdGH6vcLdOloBEYkhpuVrhvC9CrUhjPUIbyp3xY2pJfLVhqEwX
I0Yd18uzkLQMenCwY0s2qxHBY2YmtyR66mWsWBc+MjiloWR40EidTYMPt0sOjePy
oW1sCF2m7d5N1ipG2s96fZEV+T4SL6Cz43Raa5OflB5D8q93TN4xu2IsCpwdL1fM
E8jBYWA/s1Z1/TCLQKCXicuUD+lbZvjVVpwo371DOWYDoUeMbxIBYlvsi+9TaKNz
uYP0SR8WKAvFiQ2K2t02QTYaXAbaJFa1tJoXKN7Dte2V73VhyY9chNC4oJKevf/5
EDYLbEvw0xrJxtjFmdtkxRXxIOyD42dUDCYdnFAiFhNts/TqJzIGELOZ1kgUMIQ0
iq99xS77TaEV1Yx2Kg5LUxlm0bUJiSpUmJcsKVp+2R1dugxLPEBSechk2JN5oQMF
+zmSQ/xn0mDc5S1nQ1WI4EBzYsX0pc+hoqElgmLkOsXOlgiz4Qc5yK8lvSyoDLpQ
eFINJRJmKQMwX9WSUtETdcioPcdlUDbg93CF6pllM16stoI3iWppe1+LrCGMmpAd
apntMQyXXX48PHwnhcFN2J+XxhACTxTF0FYf7932u4SNK8jpFt+fBI73wKZ+bcg4
VMDd2L3Dj1uL1FPnwu49s3KBLvZmgWz2cauymy0pZWSf64yjGMSUtuwx5MCFVkhV
9x9jG9WH9jkzlIhG2BxMHTI7N7V22PQASfRbb7WE6sZJ1/FAYzeemWNN44o65XjS
us0ECkFGuTJxpsFq0ZnoMnebkgOiq/rduiI8Or207oILVBcwalJUo6UsljHdTeeL
1RWGVsYddR4DOC44EEqb7Pib5At4P6XuYY/VcdZ/t4AJtLNL3MH3xSqJEzOfZqyW
K2MWjK5jnZKPQM96T/SnJrxt9VV9zysa0YVn6v3fMMJ6JSaqfWekOSnoWJCWssdh
Aqi5UGTWkXE5D0bSqnnCE/KIwjyuSXPdAc4fmt8kvbipzlfb3nfkrD3kyzGPfo3M
jYoFzf3zSqxgvSsptrb/Yk+1UuK8obtxW2Mp1Ryyls8oDWoduCOnHNjXgNhei9rn
kWrWLxJm9FGuTnZPazHz5+yvsUYZJFZz/0dwvaa+qA1kGJrr5jwf3n2vO21whGHV
3DU1xymBJXqtLmM3aBwfEJrNs6tFYOhYRj2bRtASo14pi01A4rn4fmk0TBCDPls5
lBCMOHa92GKPhxs5Ai7+9OPIdeSAMk1vxbkIBqffbyP0WkZ39/4cxJ4oLNuX42gW
J35nYHrn8PRF3DcGd0kceXWEOcER6rLzsGJYc0z48zfThucAtW9re3kx5JEoe9k1
BK0NxOlpPxnZAno8btqf/FS9uKNELaYIKg5rG3K0zZFC/oj5zgrg8ztMi77VOPWY
1Y/tsx5z4GF0QB7fprZphuO+68egot9tY9TJ1D5++sL+qrm/YwaaS9yArUpjZui5
lu9wO6IWkKUmqcplP+imGaGfs6C3x/sr3ytDAaXMuKL1sJ/xmjx50Vmm2G30/Dxy
VQAcOOqMHYncWpCvfQMNe+D17NHV+85CeVWePFlfvwAxKmMalFeOYq/rV4pfPSpc
AufmXofhAutg/RttFHI89vUXEwiX6r9OWPZX0E4vEM+8oNQUezueop+G9AqcEcDX
LfI2Zj3pm1z4upxhi1RTHkQWodsrPhiTGvONuVQg4X0VSVXFvNc8UgChaHBg1qLj
1vuzo8mUh23HTPT15gNx+B3wM0FfoEDf+J64ci97XRBXK0bTW1DqFbK0GaHFQF1w
6WN1Y3LS/pKmNZbMp61NCcxkV/UbcTFZ5e7AasiXmhu97A2yzEXxmqTodxft2CsV
QE7wImqzPvjmY/7fWSlqLhg24afmXMUjDxHHnh7qGOri/DWk947tNc+aCCnW02Yw
yDcerKpowANdYUJQlLtMur/GcDL/qs1Fts6Jou876MWlGSdVCDVfbKrPZIDK5PBy
+gLNaHwfuutG9ImgZBFrexFqylwXgmKfG0DVj9iwUYPu0PgyaUxuctx/D0LuUO1I
wduRTbNEJpPfsFc1kJCH+OjTLpuwogBzi5p4D19Qc2fwuvTikm1mH247CTx8gVcd
tfuydxgLqsQ7gp2QyM6MWe7RQ4W/XGu5uHW7H35nR+4vp2rA9ZL7ohe1lQ+hkMrb
sY2mpcJKCVQPQJwkG/JGGaPHcSJI8jt74bbP+EVA153I1QFJ69c1yeNh03nHc85W
iGbLFImMmnE0MSkEaCTvdFF1tMsqWADeD33jCuSgnmWbaPsaVUXqAklmH5Fz0AXF
dDGTwiaAQWIpjPvqEobrxtZi1z/UQm81c8TFNIyMkkh42s6kq44LFJLh8RmboUYZ
xzytcbCbliWtYjV3fDLB3QXNK1IApkI5jEaS6snvGPzj7sRUmSVA0UAefKAgIAQG
i+l/YSk/OlIliZCCLBI7dSYNLyfF9WjamXrDnV3tazkmj6txw+UIp3F19tz/IDQ7
y5MlOLUvxdWslUfQ8DU+EwD0WHa5C3FTkGFnQY/a1cMqiJNObvQUp07nKzZ4gpcc
kfT7Ji/PNxM3ZBsx1EyrvoIzxylKh3bNpk/PKSHnhI9UPtWJjzUPa0vjfdqMJym/
VPhqSb+mU7J8bnF1yYKnbbd1Zvm4sGgFioRvm61GuCQezvwfe6dC/LLlN+qBmPbQ
aIlfqALuiVsJFy37TEHUOQU1s6RR8by2j/Ncgt3c23lUo430YKiQCHjY5rD9ohwL
riO16l8UEm0rLfBcxBA0BnMMP0BRvbM6B7rrlPxa3YmOUO0/1tqILqF2QLxmTlRL
/USWm2BhczmbzJAoPiSOumYL5EIB+oa7u/nI+Q4095qE+8A7u5ve2I7Nn0RpaX5k
ggyo4YaW3wBDEnQmEbOjJjgwS1nBokgnKKlAS5vAaKh05lYOBCfLKb67SbbYwt9y
6UXpe7XscvPYWTHDMQBZ+xONvsGaXqVdfHMIFfYa+p6Pau8EDLCenZQm1/k7YXY0
m1ir2KePquoFl8Nwb/tjbxuDt2UoGc149BMHMNDVwituohjFUBlRyIaN6Y75tsIz
UIfkjE1fySZYeMkSkCGM1NPNrzYNqUGEyPQT8+9D0eFg4n2z1SPd9La7jU22o6yl
iOKaGBKvO7GQU5V/J8eQMnjbemcZhharMvdnjqPJZfLSLWzCEi1l37caTi3l0cUz
0Qi12Hh3VBQRSg3FpmuC6SRbIASBxndPijewyJ2Ni8SM0x2tUzkij8+ziBJCYTdl
J/DR6zQh2Sucf1cv0QpR4wp0HlSXV+TcFf1uWfu7MkDrLyhlOr7BETIEbno4RVVF
Q0ixPT4ADaJ2ao8aWelnXy8bBMIXP1412TfWRJkRlflMnT4CxHweELv2kjKzhXv3
t1od7/rE0Dm4x2vWsdHONuURkEaIjC0MZkBepcJKceUWFX/a2Qz6hqBGWfigp/jW
OF+VtMRaLu0IoW4J+MUR3xny42rBFuxCTIzlhsQTZvcY3D5P0JJAz11nt9uEJzP3
0ff5QkU02lhGFnFrhZh1Oaidz/L2NgNV0GKXFUuD0w8v3JMUhJghHv7l7/g4mr/E
rIQdNJzs7ShvlE8YUSswFwHR6cIsIQ/TPF3g82JVYmez+QNM6blzDgippLUU71TE
He6ud4GkrxrXJYZbxIhYLUmXALyh91TMZsLVZT5fXK2AhOM9QJg3PFbfiydm+TLj
Wn2EhUEifLH/uU1P4m/8wwNbhrXUsXAfmSZ2AJD8kiMe+ZBmaDmscHFpvpQw7G6F
hNcEnGRgWcJuULX3DqOAe12byk33vpXzATX83Ow0tB8EWk41s3qBRHcNuSz97Dxd
8mb2zvV1toWkA8fbcEnvp+GvIPpRx7dU4Df5+a/IpwEvTLvfGBP4ZeneTQw600nt
WRpqliD/0Z/TWwtLb2Y75L+K2n+AycOugJiQ6jXPbzic4qHKpsqLucX2GgJJ1Qa6
7NvODBK0ztL3fSfAVlyQhlwUFFL3Otc4/MjcuXpKw34qmRZn07vVydpNzYYEAknp
77RtpJqpOuPN5k7Bf0xTSctboNm2inLgcz6lQFiKCCkPw2HvZOjh29CqA+zxJ/19
KolnOSTjbEHY2VB/IUKYrVHtBgrX+e3qSGwWOmE5/a5wWJOypPBbFF9cSDHWl0Oz
teg1u2yzPd2WpYTKZLySMiMAaDvArZ6y4TCa+ruQOGUweeVBODhfpV85HTSlUDHE
U22B2pK47efCAosmCrE+ONt/3qUzL39mSE0gv2SWrWrgxiAtgHrL+W2v4jAUMCZD
0xBFnTsEqYGU8h4XiWrQ7uSmt+pz+4/GLJdJsOsGu1WlLfNdIsgZvymX/QLrSqu6
1pJK3+NszLoKftIsIwJ/eF+Mkd8qMFvqeRbknuGMEN1DAZUa4KQXZL2JjSui01VC
oZ6bJk61CLPh4KSgO2DcCm2uZ+4tmLKJ8OSGmDnfKRVWqO9jC+dlpY3SkwNOwmQa
nUembAJ94qMHh92R8ao8CavTlynM/j3oqvYD5L2TSPs9ApXRvTUJYb5UNLiS96S3
CsO9J9P7A97HqSuRODOv5Cw94UphkY1u9x4haLl989Zd3KdCh88BfVH6N12DWaX2
Vn5rqssyDeoq7xEtVg+jcefFWTfZkJX+5I/mf223NiuBTkaYGA/FmTogzgX1Cqdx
tfT+LTJDAF03k89ifD3LyZ1T/a5R6TJ/hZQ62nSbihi4E177vOk3Yyjzl1URrz53
ZX9LCAeSaHmmtQA2WI7gUyEOigThslHsAIBLQ+Bv7tWKQ9LHk3/oVgZHQRw6ozw2
Ytyh/NIjS/GJ45gJsuC9YMpGvcHfhZSOoySy31LzTSAw5/cT/UFLIjLDKR85Nc9G
ETQVGOelSIc6FGcJf+atIx9agqGoDXBQZCFMncr6bXIUcSNdNM5Iq08ycilyHeTa
HvLCh3G3B3YrxTJE7KefDXAUUYxZnil/9S6dG5IPMewwixeuzm0aWBqDqzt+jrGF
QRNKacd4NLNHnuHtF9txG3pbBax1tMY0crVfRS/YZw4FWeHLsN/KyeYygxgLHroC
6KIK8FLd7J04WeQY3k4grhIoJB6j1lizmH2Xoaj6+M0iEyhyXZmPe8kkOBmoL9Tq
qPHQ0XU0pHHf88qSyEmyA04w7HRma0GERX90BT4WAloBpzIMS8AEJCLaCB7RmSpv
/sicGBKnnGkxDhBgYRtPlyfNOZLlUzyiyyUUjLq2g4FcHKSEdFYwlZJI1IQOOd0k
T+msnxiZvQEp7WP1Zviejwl6AMB+FfXr2kB9onz2xmrMKXsXX68aA7MSSEhrEAnh
BgUb3fO3X0gZ7hriu+C+u1JjrhwIExSQ/MjxBCqnX2+YWatA5h3oYtiIoAmPVUoN
jOeHIbK4tv+WS/d0MnwkEsD4I2gb+QBMF7YaSpt2whaUPZ61xahQIR4m4sqbAByx
1HzKvnapmKHXujlL+Ak8cfRjd8P85HSi1115iMgLQDEEXUH+3aP/kLvwYoXdyHaQ
Z4JntJcpehm3JKgvV2OvbXe8m8Rx4IemCAS/21D5WEf2x9AgpeKUbwap5wnTQHOD
B25X9izwOvqmVQq2vUGPaoLaIFKKtTnNQz2K+2e4t9elYbHuyNADxbqDrg5qJ2HK
4wiI1N5WxgV2LuxsX1uPNmeoXvd4TZeeIo5GXlVHOENvaF1+UTGQt9ubuDEYOTBo
uO3v+mp205khmw3aGMPONI7l9qJ397TklCy1dFd6b9L6ys0dz2ZAG8esnmOnst6x
jSVpfx1L7rlxDzhDNL0lYzO6o6JLeYLrQ5ThB5TF7/cpALXsGK/Z23nxiJ1GHIil
y84Qp9yJUy1j23RekboIrYHEdcfaK1Yf6XDmYbX11PDIG9EN8QYbumH0Ikn4Gb2P
akg5OCC8vIGWZNSc/u+NGwkuzDlvB/f3nKdhYA0Tj0N3JR2TwoxGp8m3a+bHaFfl
OWdJEZ3E/TLb2iipRu8YX0CoDBj2fEuDi6K12PWsBCqI53hst8PLISzVObLPWyEe
ZwbYZhKhV2NjNKucSbmpjQwNyFnt1/Ggi9kGmdz8aJq7ibX2pDv8C1ozPsq9bnI7
lfF0DnzxsYPouf40nuAGPsxalgbu6G8ZarZK9AnDc051lTPw7liq3VpADsyv24PV
TFFOH+Rjxu71CrcGFZREsjUHc7CjC4YBwLdYF++6nhJBFlcwAdGW5no4BxAydmQP
DHegqujIubBXVM+kQS4FlA0r7QaX6jCVDpmEho4ZeEGtBMhzBpFu37qGMBFkFao1
PyXskaNsW4i3ay+bAdMSASZ9IBXeg5iElHdn0/c+KQq+aw613C7wnWjG7hMf6+58
ZLC9qwInPfZyRd8euAv2FjD0dRucrgcufXmL20RF290wjUdcbD3dudyu7tKYKbGt
7hOB+DGiMLYjVWXiOKF28R+Xlgzdx0K1FVTXRRnh5Wiwz+bt3qMU/3PkbQ8kiwXc
Fh9bbMgJk/O8FkFUmcZdRg3vYtYOl/w86WY5yrUNObrREnq4ZBvt6lMbd6/d7BY4
X/C4Fh520IgFivOw1i1yXguRQztri36trM2ryyUVemnS4drai9RmORZyY+YYgr24
GWmLN1kdJQ9eK2Wvkn1io2nZtdT8QLuU/Y+Cod4YklZo/UNeEVKZj1D+zjUjd83m
nhnxKblFGxwDIu3zRAg+EL4h1u24ZGQbTQo1ToxCLrA1BLxjuzUso1uj6EzT7at6
obbqJmW5ncap54RT/2xLdyNcwFZoBSO44fcBfX54WYJPj8Z3jNyt+eo/Oi+vzvG2
49Mi3nyTc08hDu/j6SE2UUcPwQCgCgdOKdtolLSO3/2ILXXAwjwY0aUpVlQwHvm5
0PrtohMM8tX/8GruDr5zYSQ7MpaBFxiwn6zCX8pUYKC5xH2o4hZ5SSliaiMS1Q+t
aEmhxZp9kznCPypVRzut5i48dOucAyBFlpWpGnDHgSR8f0zRps3gIwcZdeyyskLL
Rqm7rqi6StY2jTBNDABsc5gWQxKXJWfq9vMrFVOb5deFX7yft4Y2y49F6pfsDk79
8pEqhT1qTbrZasy1d0ffOl5Q4IBZbzfP2OMrfgheDmZ6uFw3VxtogauGGQ/w6cdY
7MvuIckHOhBszItaah6qXOHS0R0WFzA5WOZQ6z3CRoTB965iz/WRL7/m4IFio3EO
oH9jtG6XVY7p8k9ViZONDfQawzumA2jjjRoh7xU+DGrmlCu5i6SE1fHLRND1xk+L
HNVB3bfQRah67M8l1e3x6MQ7sIe2ZN232Ygb5gWW1VGECG4eG+6CnqBhhwmJ3xBq
UYoMyHa5b9ISD2daXDmjyza1fXvfSKpYbPegAzJ2Z/DUacS9ImgNsN+mHj7wH2pm
D6mNIAxW4IsLASQmnx9DZfb5atTYqBEFHovGKFfBK/JnU8xhmY6yyYvNn60NkxbZ
sj9TUfzzu5mkZOq4j24LjAd/fu3KOJBek3UePxUKhAveF9Yxkma2EGG5r2n8A8Me
Uty4iiN6TmwY6VmKdHg88ljquaY3Lb/hbtrnRHLWUT6VmRyViGBd35cJY2Um6uQJ
3MzQEnkX8yfKr582MuF+ZkMzJziKsJ+exSCxw04s50MtiCI+LvxXRb7z96Qgjsti
82xaTq7sxxLKmJoUH5ZHkbzntyCWNUrbRgaJNc0Ll8WhK0cTm6ofC/eqxP0oDK5D
2nFbT+BWJ5rf7DCrLklcDWICHVTJurey20MPBxQwmb31KzJojCcv0O9d5X1yheZp
lTCSEBnIwv0hTUVzPBKJfxGTjeCTdSwe7iOpn8YulD3Wba4xe2sz/Xi0/H4sCKxa
lsFUFFVCbWcJx/W4OV5JEr2Pe3OLH2h6C1gyt14gOVCGbufh7s8K6bjWF2UYRA3W
th0fKfE39f2avcbbFWLZpstIWF8dmYt6/MrOo/SrzsFN9FgZEkkuC75Qd8cqWXT1
SnArmhilmFbah3wdZ83EkJcA5GZO2ALv6tF0rovwH0P/GU2SttJm655tGp3syJus
VV7watAdabu5WFM1NaOkuh5ofaH8PyWaWyRKaUAjnMsd1NjqlX90VPBL8q3rw9A6
wV5ZXG/00dZSd3EjRUEwI70yKLh9eT1AHJX5R0YS51H8rDq0RbdRP50e5ywNeoau
ux+tmGs3DKSuFgEh2A9SdeU+2hVvf6Ac8WJaNn+JNXwVntJX3Vb3JfYLkAIdy7sm
Igh2X70MlcAqhzIUWeKMWuCOztmiwKEPusVyR3g2PhBgUH/AI45Udyo2P3EXq7bx
Wb/x4UbHhkn7a/6BkkKHS+yI7ic0wGV2GjshbC+qOwxfbHJjH2Zpfj1fGMZV5+4p
v+ZpSJHQq6BlA8WBFuaJd+So1jojkZ0m8vMWqz0tSlG1TXRX9+EQVt4iVaGZ7vT/
LqPiHxzGB117K9zF/E3th6z0vRGp/e6HvnKZVojg9eOpEttIwIwxGNOUS5ss1JyO
I/6yvcDSKd6wB+sRoq7OcKAUqYfEZN90056h7PxUTj15cGEqxMsNOISH/7Cct1MU
0wy5StbJz6792YZo23ZZuuJFiugZwcix3cQwX+kDkdyeJiJXtX/eRSwm576yWyhu
dh8ewfaeD3WHaaQ0XpYoo99uZvyN84HYlLvMHJ8A+/RovcyrWTigw9IleqzHSVAg
grVdR0y+WRaqSUbVFho8LpOS6MoDMID0f1H39VbHuKdaGFTjQc4kQx5D4eV0rbyy
HkxJVdmn+Lz6fRd37sPGAk2QbfvWeJ2TeNa+/c1HbbzvGzVbjQbGwL8Gh6PuY9EH
F2ea/joOHM823ZdVp4TELL3Ks+4LsBbwGR6Nt/c2vm6GF9MVnlW+OlbcUPvoICEh
IxVhIqlP6ky+aQbj2hCJB4DsF2Y424kjEkb89zEN/tG5/AbhpsX2ibmVFGH5Xs/3
EAs3jrP4rwYKsCyij1JTsDoCTWj9xLTXiDJrSTMHIRtKrtbsEInaKiOGLkezOg5X
swubCchkQvrF1ljvjrC+Vl8odqg358u7C1bJ3wBZao4UcWyBUThYV7GU7ibK911F
AtKWpMLp5/Oc6u5fShj9CtUkWTZICXoshodZnsjOw77yWV6WPC+L1E1rK9ABitK8
g3gH5y7Yohu8pVkAVeDA+vat37O1CHajpBTHb2tIEIqMxx5BTNAMdHebuywrnAFu
EzXfEecmmL6tPnxx1jDaiU6XoIP6q5a3sRvhvJdRcdAmp/nOvgNcJC10xws5QR5i
T6JYjKxStP48DsxgrZLcDaWOYRxnx7ViO/uFvzUAItSjfxWOxYHLZpGLHNJRBwpW
+BXLSrQTGBD3MBNsW+7Zs5pd0ahQpjF1ek7aUAb5AlYOA42Z2cxrOFwc7jFzIwyE
0WiFfk/4SdfC+zDPMhOwdsfYL4WoFooqm0myXO7UTe4VAZEa1ezGo5u7Zm+K6aTV
BrDaGLy9Uj2tgLSnFno9YWPIGSnB8HR6w4g4/mEnrvDgoAcFxyv9StM4ADssAQgz
N5d7bp08QZLQDC3stsVoqDX8dwgILlbWAPrvEqvblgaRjoxBkM/jp2+YM81fYFfY
I+egrt8HCXL9c9o8NaIe2x1GZjis4+EUmeAZ78CGI61bPrZktDzlCKQn2PyRpMHG
D+EX0xc87b2Pm4wXVQ5ZFByg7Rs1xICUFvU6W8tAJt07bV3gY1gokRTC79JWL4mZ
SF+cyWQlaZ93klTWFkIVsw0dSc6aJo00eghr66zsTtdh07H7pOKoXwZnNuQSd0aD
Q3ocPZxKzr5pC5l6qhAKCnuldB+WOVX3Tclk6CP+qIDzld1SGA3Ha+v5uLAqztPZ
2hJrqEXfLdYsShMj+tGnPXwJ1IM59G3KKC39OIaTiQe4BZBvWclufXdSbSzUDQjb
Y2eEj4vzmx+oLlyPjTlzEyrEv7gY7uMFHHDaD2/DTxdOGKzb3js0RqFbo/L9NRFX
X2mseRJqUcIFtT3BAN8+X2MUDp+OTJLe3tAeR3DfvNKHSMM8Jq2e7GAGOz758qfR
rALNEQ8OZamz6b8nx2uQvSTpZ8CEMmPxvVEBxA1YUp188lSe4kz/bFTxyfdpewuj
OnF2NDPwE2rUcOrhlRPBIrZ6mbiNwxfW2r37QzxAwKY+dRKS0/LqBEbD6N34XJv4
i0TAxS/kfxOOPFfdu9mIcR6+vhD+LyOVp4HbHavPLCF2jK7m9edFVpOKpwWXQ0jn
dhdPssf5M3WBhFBEshpy3KBn2bmU+esCyYaP0TmQaXktqzI9XKxNwB7YcgA8X/WJ
vOiRLHqDmOxgOGhf4rs8gvHrvFWqle9EqOGmPZsKcfBY4F0oOaL9A8CLZqwzejgx
4JZ+acBvE6Fni3uFOh6mAotJcJEe5eK2g7OSwh2zFdehUt8vMYMHeMl1+Q9IMNRp
4C3XirsWrnWX8N0GTTPLIn1R5peuKyrFfhQaeoNBLh9IhvKPEnvhj5BeCJrUF6MA
qy+vLRwA0mM6D38qmyoL6khntqH2U6h4nXdgFacui13EP+BEg3X97IZRJisxqsHY
Sj/rIV8ZJZWoIoTZvve0jDQsVx9X0oHKXTNE16DfT/s76DhY6Egqo651jrn1+0L0
jKxn0aPy2rr+NhD3LUCj2inU2vuk3s8YapxDDmjD7dEyJym9UqHVPdVO/EYSjoNm
WrhylcHGn6S5pK2rc/9yggOjLBflS8PkBajEI+LjNeqmcwdHIt7Z2Q47QEs0LjZq
dglGBsdxt12uIlP7IvAYtIooN2/tqV/5kHTYgDJFDTA2Uas7aIJPS9hv3KKhubpH
Kqya1fyt3XfPXPMvwIwRIzu8GAsY/il6h+oQK32w6uGRFwmdWLOvk+31I/kNwUOr
m0bxwA8bDqU2qI+4YtUXIBi6ydkhkIGAfV46g6TSvkGygDZc9gq9LQWwQHLxet6U
a4RPLn7OnmK9SyU5lngI8ERlDveX/ERi6Gk63u7zmugJ+QC+9wqTVLamGhETrBO9
WxlOmVWM6H7dc7VosE3EkJy24WNHk2RGGXi1RHOOmt8ptHosK7T01rm9tvAeFqV8
+mjlv4aV1SXY9psAg0pUqtDm2mFnoh4HBnvUmpdF7hQZoGWzZHuv7vEwJB9n5K5G
74XNSWolKuZI73hgGIqs5oo3ue7Et350BfOWvOcQ260KnN1QycWueE/1KA1r40oV
pAZOy+wpJj3cFB6vLcb5T3Gp6BJ6YAO3tEMH6h5RWxTcSnENmxUe5EeYrxTc8Qn5
vR/TmTcxl72gTzbERwwV7RSmohR2mHoFe2QLMJ5JQMMSNpwbsqFSKu7187tA21dx
ceEpcXaAGXLs/waoWcZoO5FoSEsULD1imzZocGAETC/K+J6mJEjYZ62ra2r27YR8
e+0CqAPf0IGoSBhT0Gk0i1Ng7J6yDpPMKkYxge9x4BxzXbXqUygFL/2kclmu1sez
+9FHbPK2Z2PF5R/NQSCFQQpQ1Us7UQj8N+e5CGyxpQ598piLvrrsUaJtXjF2jEE6
7fOaIOCIEV+zVttHft0iEeQ5e1Ar2rukRKufZ3Qq7eMT34IF7Cs+bvATR0dTgbzs
DhkcJZfGfI8k9T/3L9eIMx+ts75stkb3tcUIdNUvhV1WLmWLQhLsNZFZEqslcm3B
f3+RcY2Q8S6rfkWCLnEtYyHQh7VBS3fFG/jSQdG6XqrfbtIWphzuHK9WOgTZ2JA0
RO1/pX6Lsu7zHDfFDaj/gJa4SUZe/WaQa5pHZviFOc6AedC/eL4q9g5j/aD2NEKR
HGZ30QZyymyq6iIk2mlCWz6oj39IRCX88Are0vB7JsSHJzojITCf9sZbGIurJJtQ
mxOp2owb71SDo9BTs4aCUc3DdXgo5I6fMbpsXSODPWNVT999iPXe2tJMMBKEagm9
oIC8oHKoUu+U/EtVd8JTHhpQ6ITqrbC0zRNrNag39wzk7NSYw+/fFqdLYt1y2zPt
Esm8kOHF3xA8DCFpO0toCyLlsPyu/ydPckxP/zFWdcsXDwejEfmO8N92OzvSyLeV
6sxrhWMkVd4XDgoAMVC3DB9BPo1IYbgKajlB63a2J4qAxKIGPFBjZyHs0+y8L9xt
WlsLU/ETQcl+HfnF53R/3G0+K8Mujiy3NN0g5t7US6PeXjVxlS1JTQhUuysF4poz
/f04EhckKF5sRZ+cHt/+Q7p9zJ2+IeD1G9Qn/j9ns91mzcNWKloglQCTp/KdCrlc
owCqjjrGAYWMDr/bq/v0u1D+lRaZmIJ7K5KNuClSgrNjHQAyNAlqQyfu8AYSJioZ
vClaoIVb8/DQd0FoM50M6mcmwVGj85sSo08KeZAcW6GwbsHTsX/Mul13qW5Yuusk
1cntm0HYV0w6UllNvLZofOuO4AD+TIW1VxNZAhX6196VtXsqQNnWWDl3VuNDBAmt
kSbtfDxAioJcENQttD+Nv9SddjzA4YVkZ7dCx4DPslvXancbIQlKBPjohnAxJB3b
CzcXWnhybyExBfdYGlgJSzlEkxR38C9LScPpeoPZatJDysO2cOObp5GfAeQhZBxa
uzYdnIkcYHZCrq30Uu5s6mADj+qWdyfnUctdwxvlhvB43HLOQP/T8gfNgArwTAVx
I9A9+sn64u6a60ot7p1mo7axa01apOC3bvBaVZA4NuTIN4GcSavN9orEWbk+q7m5
cLDGyO6XLM33SWQuL1nT4VWtmc0S54qv1YATYW8v8qKQgV/RfHP8NfZi2onCTf9e
gqUKaWdOu4/5j0waFW4gxMMjdV+/x9gyUK6o5rl6mkn/P0c4bJIkLZwX8Nh8iZdd
nQnpzO4wYuMSlXxkNkwrwaM75e0vvkOX5z5NAfoXS8AkqdlUefKEnaLExqboeTRU
/e8+9Z6S4dsxIwlLgaGac8bv0xhxPK9ZDpAqG1HKd5eTg6yc+M8vP+7qEFJU9JpJ
kX+H22514dgoy6pB9K2znqqrOVwqBYj60dMZa+JnjZwKQd09YrfdWi8LvVZ6p/2j
kIKV3jedKjehNpCHTfvmBbZZ/p1jgW8GY/4c2gPeO7+S9Ywgj1wkXz+Zg+2sQ47n
M6p6+a9k/5tyBGVzCsjRAlrntyyr7Y7TMHf51X8wWhCc1dWtImJMAPnqGXgGNvkw
5JFEcdN/6BEt2JqkHlNZnlcH2Rg7ym117J/RI9wfzmE8c3qThRBeSAuPB90sXRXG
OaKUON+VVEl7cQuUXsrEn7B63IFUzc75BB/hcCG65DCADH98aZpEMboLMwg26jjM
QroB8yFWBqWVmx4U8DciH1LbFTvLKNiaQPxHlwQTEilSy7iGSiIrp8l7mD5TK4W8
LYvJqTqOI4Uz278uPPNQZ/mX9a9zh0SzSL0zLhLRf+MxJBHWYotLKZ5GiopyjIs6
56VSr4Xl44EY2Bq5DLp5m3jVbllY1jGoxhp3TJsC2Q1AqqBKOU787hGcdyKe1Oah
J5uIeDvE9CFQoijAjY2K3as3KWgoolftDmLZOe+PNLO28zyOcEoL3YAtHV+ilGzq
eGPF7nJymG6lvlp1VBAQEzuGnffxWG6kd6mp2rGvSP2Wl2VsRxUkBaL+hQgLccKK
Dj6t+aVOQSNuZuErKVTKdLiDWKEzNJBcOavll6ry2cNBjDG/4+vXMS8Lyr8DtYX4
zAnGcAycaY1fjHMtCLHwCft+z6Uee6mGmmW8+1ZU7Brl6R8uGEmgixLhYesLGDCT
Cf/G9WHDX++eV0St/9oKlxs369KZID7FJfPSBR18zo6idl0mpoIVdkYQrETLgz3B
Rh6pkecDiKoPxpsGGjbIKgMBSc81qit/y7q8v7PhS8E7TjXTiTT3N5uPxfpp7Wwa
+gpUl7f/7s3KGirKyzGL/ON8xJStTbUqYnPX0vwNpdXaXQBHdRQbgbTCoiqJTslp
xRtA2dOSG+OjtoedA20wj4HlA2zMx+q24Xcn+m7xnbbGNmC5kIMRSdENFiRpMkCJ
tiSgS3r9M6ebGSM8c0BJTN1/T9ZQ0xAtfvt4sFTblmtoE+h9aZdWppfreikERypC
ZZUXkmywX3abCLj34fXAK6ezPUNaNN2IcWGHBc9ZCMsWwb6gw0GFQq5VyavNa16W
wJAgo/XoFW4pmZPEwQm000V2F1K/fkkcl8UgjK/gdGwPXA7AOIgoc8j2XTrVGtGz
nUCkU84sraE83N5Yy6osfG1K7niygphqhUkjXgBIKXt++l5v17rFN0hzFN4u5GXn
UrhYyk0t59w0w+UcbF+eOHeG4E5t92c5Kehtabc29XbUq1bGARcOa3S8SYVwQKpP
xArUxtJr1MgUwxQZ42Q1Om/mG728KlqOXti5sz82iDWoJdIAg9wa5yEVeu5E0fMd
lExGVnO7r2xz0qjwcjhz1PAD84OwmH2uhjB6GOrylsJ7diQv49KnYELizcPdLnQL
Tryoo0T0X6swaUv/UjFeISpr7IjO3V2QzyvzARTmnNr0bhbj95FQtL4k+RHOCRGg
LmYKt0ebevdQUaEYey3s/YmRDUra3BCleRI79Yon2hVUMJBVelRNYf4rdm/zVIRf
y13VevXJOecJfnGjf1grXDrqeDX8T7gGxjunIDOtpUgOaQO9/DFdWZGlqOhr67Ww
9IdX8IMaPRI2V0K13KxdD/XYDPQ9cRlmOnEe7lYZpdj77Cu5Kwlk8ONtZlh1Q1Qk
4WWo23iIt8pYrLm6/sybiUdx8+LMvkDtr3pAz+ZM64+rVQmGzBVLpktoYNz/EqhO
tLDXXBsSWnFrCKkowU8ddWm70C16ghH1ZsQYT8PyLOondH4lp9A4Hfn7vb/aGKQP
XgdDiUd+lgCBYGT9y0aDey2NU4ooSLLtjmdbF6lazIDiczR357KyVrITEh4ldeYZ
cu0XdUiUG+bgj9yw5hG9d/0wxOk/e2XSn2f7BcVFNF++n2yW/QhwS2oe3F7BsnxU
WhEPSK0jkh+Aq9bIE9NOwSeJAQZc3LZyaLV7kARawTDjXzFxtfAErm/SOYiMuqgR
oBtI2D6cyVYl9XA/8+ni57pbO5V5B6i9e+vKTAJ7ke0lBH6lKi4jGNm3Wwh3kEXk
hLmPI0V03Nf08Gz5TfmxdmAHyJ7H2788e2D0sEQPMVVAygnrTf8Ew/5KKbfE76yK
nJYe5dQOClYIBmLTuNiRoT+WjVVDu3J72bxY/5AWdvlu0HQExqwl76JdAZt3FHVb
zCDKzC00DxkEhWZgspT0uH00UdXme74Hr+8wsiTxAIxJMmjGYCJG7YQhLjP4cYYN
I/dzBgLBaot/3zMPevtfEJjGzPbcEyJBGEixfC7FcoE1y9+Qs69gtfz5qtdLvxv4
0r00YDshEz3MoFydu0G90i7k+OKa9LhtyoHO5J+LLem7/tALKG2und7ShE8ZBuXL
OurAbPr99Cnua4PdSxhVSjBThaPb4jZ5NYJaxJvYGIZAxcIFSMoZLBqReDJdnuGe
DDLr77sPzk0L1mjrjDoUN1Aliym8OmsNC1963DEwh/QDg0bDcEMNc2PqNkZKRzdX
LbGJaqPjlDoZKyLVmhCXZ8/qga3cpmq41KLPQLiY3ltyyaFhFisSVDGsJyrnVDPC
zKt8rGojf1ABi78LOYA2zFCnxOK9GdhbU91DCzPHwFXiCYlCYG8cR/NAvL49oPiH
z3N7byzGT/dpobWQVgdJML8f1DCAK3KAXmya2aQgwinIgXjr72ohJUT7tVQYlLlM
bE/uMl/cgGc5uFl0rpa/lfCBCkVdOT0f//qkuEECKWwXBuIZABX+2l+WugnvHUyr
ojJZJjQQzJB91MzAj5YwOtAsOk5p1FQ/gPZX4aeQdRUVwHRsS5polLyfhRJnih42
XUbdJoDh3A6ZgV9noe1XPP6oIbd+KqhT+RnKU8oAh+aNHhE+RxxzGfyTd35XWMWk
sraqvibE3tuCyz9eZhx3zUF1LDLKhyA+FsZqjv0B2DNzDNQblHZCxqHtKuSEIJtJ
leNcS2PQdDNwZ3v3fngUdTum8ZeyhrWHLDKXVRt10PVdVcJGo/Vr/m7Ur+mLnUoJ
Zi5X4PPdVNT++tILVKh/50zBga0jekvT9v2qRRTAMs0OzpqOhSjXP1ez1HxKF3Wz
8GvMmzBcygaOVVNfC62tlfwIPWB8H0hr3gwPOgLcyKFu9ImMcTm/QBvCW/jvyCFz
6zLyLWRA36vq+AC5Idbiga+9tq/AKKn1miklbV7Bpc5g+Qg2a637YIzE9nk3Tw3g
Sx6Wzzbju9QZ5qgumikYOIy5Q0pa/6n6/PY+rjJQGyBjNbUwmAy9eN4jQmcHJdKG
sDkI0U1H0gjedepABbQZwhiy8ZEaiBihPoOuRpq6lPsv1iHvl7KMtG9oGjW1qpgI
qDQHFqWiXvOMK3qagt3ZDM0jxnnaPuUQ8rzFYf3mat5hdO7s+kxnTyUdKTx6NAuq
IulpcZsYb3OEk3U2bVNBjLih8Ks87UUWyYzDL4w8ecGyWXvmvKnzqZfGHyH5dx+H
ukhJQan1+vVBuewqAW1baw71RSjdqmHgqYQSYzQ/bYRriE8FBor9Wpti6KH4M43U
FHbe02X2qZ/RsBuWcpjuHwjinzQeYLtKaMTflt7pmaMxeQiW5Lxr6YSii5d8IeJY
7z9uDbUaJ29IpvU4o+l/fjhUFFFnuRaJNKyMEhPXdlJl5kc/u5kJjT9INkgOVQ6n
VPZ+pnC2vOtdXgsO7QIqvNDrMDbTnw99fecnb5KOmmnIG0CKXjH3GVAqAmZ+5w7D
DS7FtM1gLv/Nv/KgEwqGVTcqXbgdP/hU4A0lOcN3a/kkGtYONtI+AfA7wEwjqxR9
fkKeG8lZJ4OvppUH1UAuT48jAtV/Z7+TH+79/e0qHDrwoLcdteGSxMCqLdeI5N7x
/yHqru8i19zigbzvV0CsiEgAOE/9saU2jDYKAU77744Mvr8he/Gkj9KYg53HFvPz
7NIeaLdwV6i2hqbHSnX2MBkRqNRS1+Ho0RMoiqqjz6UOX3XUoTnRBn2QCPwkjl7L
iUuGEX1W3t5hNJ7brJxRf+5/K4JyGOIXYc2b8WCqzR7/TThpSERSSErDQQE3iZk9
TGH/UhUeERnqUaX0m8NVzxoWWyBWvXD7qLCZUlPjUSOHF40Rq/lsNn/QddZlSSUj
z51HTRRejCzQ0hKllNzwjq9GGdDuRRwxXqIIIYkcg1P1HSVV/3oNPnwUuf8qBZdW
pCjMJ47OHjVMIBKguv7zFQ6Smpyyz6CBG/gCXs1DtpGhcbM/MxjC2XL0MUBel65v
gduUA1cwk6FySB6M/avGBRxJg+twq5Uz9wjzAjzonUp1uUMmhW4S5E4fjbX+XdCA
mzzx9+Kx6IWQHqBTOu4sMt4Ww1C+pINZPrWzPWiTju7ZVZvKciIejiX8Tuwb2LcC
hjShwKEd9sAqdqn6Y/dBRnvU7mtAwzFXrZLXmjJgjmC/FryxXNRGWYjqjVrjW2GO
rwEYAaoEUY7Lh+/WUgZXglVZgu4d2T1145aTNJgKJF56rL95HWL5gFlcLRcYReV8
cIlgz2n7M+WXI3Bow5LjWJgcWdnLy5r7fhbakx2UrS0kYFs+O2nll30DpA8qhRNo
a3lbWdfOnEKF42lF7iWoxCRmJWw0ROoH4pkx1CyNAPqgZGlmMN0Rdj4xdIe4KHa0
kke/0dsu+uPny4I0qGNS+JkH71FUVL5qACsWjacdnp751S61zgjIFHojcpdxTO57
fIH7kYN6nOzg433TOiCWrtrO1MXJYZ43OFD66xucOcb3wmgJQAj5h/kctNx9Opm7
mkHyJjMloboXZTz1frZiIRs1T4ht70R92rheJxnGvrHIJ7UjvxqMbQMMpyg0hXbf
XEAZEEhh63d6z1jxoJNaFeZpiQqXqqZAMRGYUZ/NJUHMIRF/BGDqwiTbzHT3djCN
JZEFi0Kn+pMuSGnU3poftF7v7mUwmCzqYe1LSADdiLq9ufJL6wTswb2hsZsJD7Cg
jkDevYPPBFRFfRPmBpQoEFPByH5rgy0xl5gYNAfcqCpGWs8O7jnwyvBQMQA3Bg2T
EMe3S5Hm7NnmpEmjMo8x6b9Orme+17beSK3ntSXXS8FnHvtf6DVrSqUw3uzcbd9u
2diVfY8RlKOjCjlMe5aa2hFyzC2RfDQbRkG2Spnugwi5KIDJpv0ckqICgsrwgxZI
IgLI0RcWmaRTaCr4++c/mE5SwIX43MP0clXtLvUJxvrqjAjj8vhnN+0OezN7J5cY
LIw4VYjJemzqJk2ALW4JfWI8XRTxLf/v8FT1kOQH957Lp5LDkH5F8m8J2vtkKnIB
BwpGyRQP6MtDAvla0P6v8oVLo5Pcl7PEp4Pr2RyWZtrN8YbnTBu84IWc0JCh764h
50pmkvnCTq4kVBOvpCPmaAMH4tA3krBhU9H6QKSPbj9Rh3Yey8st3Ix4MC56yL7x
hveXO9bXWWMMh7Rp9k/aFcFU2ckVHB/E5ZTSr9A3qg/goFjkKju4jh7+kHIMQGON
njpgKIYfK0hvIYai7UuOGtdW+AbA4k/KO7h2Swy9prCQIvAvl61368nldbIIhgE1
jCPEjhcZ9fwFPCR3xbrRb6hvGYKJ69AXvIYTxCL5xfPVJh4c4f8EHoARJs87Ovxx
OdHnEoMMZSlXd6R4B+wfCJlIN6P/O5bLR2ZaYGEGRvOAvAAx4XNjwK2BrAtSAN1H
y78NmjB8dwrViCr+nZ7F8NTobPoLHbHrwY7VLoRn+AVXEwpInVFCPLjorBNsjP8I
4XgmJP9w0hAJYT7d7LVVWHryIoWPU9pWV0/R5/VUQyrdyuQ/1BHe4Edq8by5TbSt
Z1yRyCDRtu5F1cKgJJFDw52F8bEiCLOqz4NAQ4TMQ8j0W0NycrMqzAs+5Ae6JTBZ
77iT05UG4SGurSCohu+iKIvHqtznnIcAyVBpN++SE/cjnYxCVPE+Ed6Kzfyo1atT
2VVco3xHTRoi4+y9zcvHqq9r8mlrQDltj6PJYXDzU4ydCB/9XeAgJWQUSRAPLEP9
W3c8CF9mXgQyn6n9GWkl9UsR2xOIuQWELnBM75GF4pQhPZUk6p/waA2A2Aq01oVU
ShyT1cclWLTySjquCYSsB3WvAdWPGs7x7su8TLggkCb92SrZV3Lvv2pc1g7zsrOk
ExJpTT+IxjnwRrj3w+vQ+RID5qsApVj7VgOe0uAPoMy2gdkuFs2cACuMr7zMe0Q/
s+AmWwLaHxAXWL3zDM0EOeL8+1XWTeXf2GSynjQfFjAVeC/aiXJgrQKleaKQ8e5Z
il48MRzKU7F+EMGJOVgYrXUyvPV8MiPGDxjOTFHUvKimchjTEQq79V5jPoFhL4Aw
PakV9I3pqxAd4cWya99DyV6hLyFtb7fxu37n1zwPjAM4QJbFd0zM4R8e7RMwq4tp
3iitdudr7jhOAOn95GBQNsj1Xnvfft0GOOsDWtTKW6R0qAwzpaGncCHv+RpGZQnq
BfvJK7sdRVU85baNYmTOe3SrcEgRvKWTe+wOq3sUmKuzIXLlBVvgGpC2n3ZfT6ti
dK5W3i5JNN/U1i991hcX3i3wj4na2eMygNcyEV8ISjDdCIJ8hN1cPBFuVxC1OCZZ
EFc401hPz3rZ0YsMz6kdVua1DpXCV/SPCaT9dYHkwga+5k46Ai6VvjS2f2qxyXbI
iOW+MS2Lh3qou3NBT9s0fYBXrl8e1UPF73S5qn/7c9QQ45YKMcJiYwq4pMWctt2O
RpjaeBSumw4Fmn7NIomdex9JD9AiAWJqpQpVm9SnG623HcwAv+XmBuQ+nEcqRsol
/PI2irWrRq7yYBdF7Jz0fi7SZlv4Tm1b3cxY1r2vxfsZ3r4OFttwxGlaWr64eRf4
Jc6CbsBMs6njQJ5UxuyJcZ86HQKzwymYYzGYbWW/bM8cg/N9siKcCN/Q4h4VDOAj
S9DHKF8GCJ1mtaBd21oUrZBOf9yTmZ7tzw++EviVW2ZYzIzR3i7NtANH52PFphvA
jZgxUiARtSw+p1L16LYDOVCWhsTyrEw25yRQNy/zAP5TnMFZMqzMHcs/SkQTyl57
/gV4rHnlqwb8AMVP/RCTTgjsCXKQjyzVl+PvjZHhns5NjW61l97FS2creq3T6jkm
q49dti0+H8TatFpg3ZnVhGaCZjrBRKboV/51F9S8uvvG+T/sN2KJ5zH1bP5K/hq4
7WETh8jgKqBHILGVKgUahNebMUawCbnjdVtnA0P6TwJNMtUAVSpvMx6ffAC+GZqz
ZLvgOZteRw6g22KMxzP3OCinguPZ3cjKiNJIssDN1DhKJEyeFi508gm7bJF8GvCv
I7dqWtY+pYTRNXG2qKLy8d/R2ondXk2GH4I+tWAQdEOvc0YOV1nkjbPSpduRiQ72
4Lr+0U6gTiHC61+NxUQyfHo4erLeeEg9NEzepD+Is0U1ehwZ2HJCz9y/uJ/n4sFi
jDInXloqK7NFRe6kG7/UxEfGmutfRKybSt6EIVII+B+NE4O9nKaTl8iz1nQ0Y011
adtTllz5fpT57JtwHpMCavDHlx7XPJCUVJADUX+IIDovSiC/dv7qiVHbP6Rkt5oZ
zjE9tGy3i7txept4nqJpAOcztCAdxMXm1c22EA3vQ2XvJ2gZlhbc3FiGE9WAngdf
biGTf5fp8yjg7kojlFw/Wd9U8NpHkareiTnKFKTmdYFaBI+9k1TgTwu52ecRZRri
Z7JnIrcQHyZ8+irSDFbLsPVOPvubXnQodwo9/ilHEi6JT09/FxofI7SFAWxmglGW
Y1/ILx2phGJPgAlurfONyDqfTfw73dkriN5KAC6hPU0ZP+youN2KPNvsaOX26ebr
UXUYscA5+h5dRok+NKQkW7aGck5npcyO2Gv0/9iiiJmkAROk5iWy0NaSo4fK6WYJ
Qm4LOvHilpLYdDEr6UcJMa0v1AuxpBUDAc0kCcJIRXe8HhhCWYihAFG5hGCWuH50
UgOeKOYLOWTWt8Nu8fJEj6VooJjADXQ7UQ+1gihi27LA3Ujl0bSTWIIbHLuEUxYk
Xxf3z4TBAsFvfKy9nK8qnebB0a1iqY+jZd4uhDgELmDldmvrywVOjT+zs90gqIrg
nNvsWLJFDqIldqjrTvNo+Ub2QTtC3+lSM3NtcjROg+wor5AmnGCscVvkdZinS49P
tIJmDuTR+nMyRsYzyldPKL46Nb4gmDG3Ud+oVNdZUZLoh1kvju2n0p1EhL0F0AW4
bwwVG6REeatxc7y489BK9incRJb9I+BI1Jb/BOQ7ypki+FpLnAdu3V2pvMj0nFth
WcoDuNxx+9DrcL3Ltyrjd08RKHJZe3Xxs/dOcWVdWsE/qykW1kkMkh4PLZ9GYBEt
nNQZ6ahaPb4FbRfZGjTk6APlg4PD4HcxTqZuvFE+d0mNt59d4X5lndO0Mt3nyW0C
MBqFctCBG5Vurczy9ICenACaiqpXGN6SAlMTGnKKT5vLG6t0rY0xYe7+ZbPQEoGX
gSDR0fgUnmkYRxqHJzeyT+VfVE0sXBmPdGNNj0TcU0McQF0Fb5WxObnAbBVFJQsr
U9522eUf40IA7rsLTlg8W8Zrs/ejVX7a3b1hvkg2Q/bpWDn/SMnB9oOoSfL4oIlK
fMNdi44s4N2NqiAgGwKCNEjXC+kMGrZTKT+SNPUnj/QAABDJLsEI9t+H1/AcyoAM
6HfOftcI2qWDKhmgDuHTpWZF/QVPuZxaVplp3AiCtJUCAtRwq2QgNPDgKRpLNRBq
njbD9whNBIt5BXoMi8yDxIZ4RCOM5v8EseQ4PLxdrYlWnF39YHmvHdetPlpK7csw
YeptdakalVfNxwcsRwTaPe60WyeP+M7N3DSOaEp4TBZMUE7Fg89W6oBkvZiVtnVk
KyDw4Mj92lqxETs7/uhH+6HqC/De7+ut+AQpRvO9eGSIel6pUslHnvlm2ZLyHD2t
J57QdXaY59AGnCirZUHTha5t8bFoSPgTuV6kktcPwhib8ZoYYsywoUjZT9G6LZDQ
a8O+ShuKwZ59dWv9aLN9SkyjErD90MbJ6+7eK7XYAW14zVsBYrdmye4gsXmu8wa+
UoyL0QjdgaDcL7yEiCTSMyGrst6XA0xhEwM4USAUB9tpYCOn4V30qxqnnFSR0ib/
pLnLQw5BB0oM96Hk06gRfTG0z0VEaUWR+CyS2dyACJ6rZY9tXhM5qfUbKnNnCbZp
Q9X/gTaZb9OuGqM43vqtecXB/WtxcsuPy9eJf5k5LkkTKrkMAt0fWw2gHZw9+tcw
ssYSUUGqMlpcjxhXcaoJu6fFeTVm+tB1zmjNKwK4HS/ormm8RTLVxBMuEOSz5WH7
/ImG48E6VG8ufpmzNcOo80a1wp3K1Mmlah/G2nQ3p173FuRW1A9AWDyZS3dRCLba
XMsUoA/RhBkC37UAHWdT0xmM2iUjZof8gePaWaIEeaUnHr3JtWHH/o7WZJHkigIL
q7wFos/OQUd5KqfNk1GkuAxRhxks9FOl6vVLRVtstOYAUUJHmv5k09Lp1QqKLeG0
VyDPdoGpJoawe65u43c+EHvt6mcbu1MsZ/R8ADt1cyJ+Yr7s4IOvfYeEs/upDnH1
XYHxYn+36hbdgtO3XL92doImaWNlGgdgrb7ioWVDDn7ttveA17jgT9IpesbQZvZI
Y5TbPuUBFYtgDwrX/SsWH86/tg1IvT+WG/eoBOtfQBV/BEB87f07ILqhh+X41M9b
MgDmu2qnTHQdetwA0SH4pi7ONuaD+vfxtXvb5ohXTeg8655szSC9NPymckRQnkkv
xDI7jBE7d0tlC3Z4wldqOCX3iOsbXNt65lgSFzbcu/mCSkA+W69qCEdJdYmnvdsW
ZT6YfgBMMZQL4zXSVInd8on11cf9vFJP+tgwG4XktqvX0y6/MjOnZHUhChmZTH6I
4+vheUjd13WTamUeIh7Um9/xACha6BkHRLH0YKuXksJO2zEtxIJBjyq9/igM8HgW
piGX3stjVSmZ6toaKOk6lIEBcybyKCr7cj16c5rRuKNRGioBcQhduqqkNSyyJn7q
VvZpcxsxbzasCd9sdXBH2PMapJADhm/JikW9nE8jnlbtVOFRyDVdZyL4LZuTEI75
Tdjix+sDwV5yGNPRC18xgmFBYDnr3TVZ422fDK31vpZIE19HhBTvLYCFiEpo77sl
618tHRV+nmFg+hI0Eu9AzmmdhsrwccLQeUXoUvKkc+XpDrar5M+zWmwdXt3R+q0I
pt4BJdf6wwKbjrb7G4g4b+onepTrwN0FwxX8JVld0rOErV/E69fEKSRqR5BwYFEC
Sh00tUV+fWB4p89xtMVo/dV8FR7tPYju/Og+vox6b8Zj8ixi6IyyvRG5AtnvV9Vs
FxNeXG4UCE8JHFmYzj1QAVfHhajkCwc9Muz3jFAmxtmODuTSsqEnP/pxCwGqIEEF
be0LQHhZoI0qMtrnDi3L4yjVUffxnQsXr/VSDp0rJNZ4m0E807/VxRgtYYAOvzei
rSreDXfZ5I8chwc4sfl2FqriQlw5qH1RhKyEUdpnXvdJAdcq03Q6RG29YF1s5+51
hxlaZ7LmxDji27wnEW/qcX0/1KzDV5FX8iHGul9XKQ0lxEgUkK8QNpJEa4lXr8HV
cbMGCxtkJk0WeMC5sMWZzz/ZtFgJZjqoVj0B5hy1Osq637iuuKg9yeuF1QnWtMET
2icSg7CSkhfx8ReV3IB1RQdiMznDHFbc3g6RZ6tFUAsskMUnLrW1SQCssa7tyMU8
tZKWwbsbXrBgnGK7i0BpnIMVSY5rNiU4K3Sf7M8/XoUdNMLSN0CzWqMTV+zhLXM/
A1fnUp8NCaW1vK+3K3ffiTaRd5pLFg1X1HtWk8cxP/CmxFdf60E8VXojMHDEKxEZ
xlwsE2MlCSaFrPa0scVLah1aMPRVEbNeBiMOHTwDJwjWMW1Kml4jMv9LSlZzha3N
Lu1fTGbggyCnoz8Zytve4kKNGwtVse1wSloMJPqHF/7mH5b6I6pGHQQAO29gzv/Z
MSigpFLRIc/9QuSKk28Q4+f3W6T3xpjZ/jAOZVbEr/KVn1kKyRsoPo/yPIkb83Ia
YnrlWt1rhalBIyEb4fB7MCCQMaNQc0d3MHXTJrLSPyiapiKaNnjOY+Ux+bHgLr5O
STXX2Pgd8yYeckLeWBWdWj+kKF7oMO7J+I1mXa9d9ms/k/K57iXZpnDKQPJAQxsc
mh3Pw9YnTXGI0nONmUPhCXRSVAsuBAnQ/mOJ63nZdxpGI/N0ajnuvIsDZL/hZT3s
+BSvvcZsPIA3zE9tQk4ylD+E2Cpxl9BNwMy3hCkDlrhVK01enNlH1hrgOmTAp/pI
xp/nIG3m7kMg+/jAGUYRRGAdEL5UAGZOgiWe3ZjFzdfquF9wwL0J64vbeCCgJHZS
XmUCb8qkZuPMB95KkffwOLZP2WbqGOMVH5DNYcwLM64fjhlRkh/uFIdqK98LFBb6
Nvpc13W35CjJubmJnzR4Oer+OkexrP4YdsMO+PkxnHHq2ZEWIyquyEVklI3hyMSD
+1yx6SpSaTNFaMRe+97l94SkjgFt7l0aFr+5wFKOv6Vg6IeY2C4OhqB53jf7k8xp
frDUD6OZIlqRhDAk3IizsNgPs0wgOyy36Ym7LE0UIVoOVANEa7sfEnRCkS1Mjm5P
J9yhoFfKLOjC1cb6wjEAgx0agFPTH4DlpzyYZTSoltZ3NEdGLqIAfy+BHFw+0Cem
xQkKzt079BLJIJnaDGqF8WH6cg3Kq/RG9DqSwHFa3knnxZairL/wWHBU01bELD8c
pVDal44W2ZnL6AOM7iaqvJ5o6Yicq2I+JXue+fffMKgk+8N8BfYIhOCqaHk+jQ+L
pESc0xaVibjDRUqR9SMb+jp5cs0xCJ8KtV7TsJnoERdH5CLbYFpcwrAhNF+aOXEN
Gh5hmYRJGXIdLeQ4aoFNPztPlPJixIjNVn1ZWyow+7FYXcp/PdDEpmS9rsHevlVD
kQNGI1aNcyo4AyH8sQiOjyonPiexNS1wuclyriBuZxtzDj2e4RCaLDai7+Kq5JDu
7nQ7JsuIk/UTu7SaGdl+HkIf6jOH7Exhw+0zimNOKUFOLTt6ZTezSMehFTRghXH8
9FvP/v80MiQ5KPPWvPdsDF2AFDluTuHT0Q/ffAB8pEqKwdD3xmyX4Sutv3qS2I/r
vOwbtm+t9X/U3sgEjOUMogLPWUetrdfd57JZSaBjcsBdsHzyfHPN+9D+7/DoNmBg
kpckfbvFT3GjAaJIiuoJl/mGUZJ6ZqK3gHIoPL/NW36nVlzdPoRIwDZdWvRDvMK0
EsF+DqYJGdIv/ngJ0FknGpyk/EJKO7gilIvAMk1Jeg4iuoEoaWSJUBjRCU8NC0gY
CcGUBHq4Fslt9exJR/irbTPAj3qmE3RvpRujg5Daf7Chd4qyrqVnNP5vt9oOq3Hv
kEjpxfP23jn9kZALbmFnaZV7LOT61Q6hheyRKqXlY/PY9xr7o+SGgV5pzh34jwEc
ZHeFpPXhkXYOq1MHNNraNcXEyalWDv7QknVJuSKCKFEPzUcAdotXS2VDhXopysrC
3/zphpsaLHDQTyfTzjSOZqTHig3KcqODe6EPx/mbl0z7La0R663/bkpy3ZVK8Bqv
RQwAYQvO/xEAylFnWduoVX2c2dxbZJplqGCRTllrE71adT7PeJOD5MOBwIYpS0dH
urX5m0AxOmzot/6PzuJT4Fn4GSg1mHQEM92U/xbdJJgNg9ryx9JPf4vABDC0SRKd
yeZ8HcXld726WxFw9Xo3XbfdNUdxs3r2mvZmfzLKecPheHXi6j9AvKPURNlPV1b5
KpG/NtVl4lDkPE8JKsoUuVuyRyjReH1Gm9/7CIAaClviIB3y7WuK/qj8sSvO9onm
rPy9bwCDZ0CGW3nWuJzw03vAajthlnN4hoY9I1CggAhwKJYKzanUFeEG/N2o/Txd
rDsWDbSv1c7qfAf4deQwvYhNlcioEDU1TD5k4EH6NIx6ceKcIPcCT3MIeaDd6dRg
CjFGzknxNgrlInOQXFFm7ovBLA9uMNfPCfV1G+Q5OtonKEkMZM+Aay80/I7oQK5a
4GascScfyiyp55j6cSk5YYw2Uykoyg9ZKlvgelvfNEsVM8Z1Vw+0klRl/tw4LzTC
fcmbzB0B3QWp6AqpqiN2kf8w7jqZ3T3bK9lLgzIVUKkikkiLz0xlDu/aFoJo0Kme
3yxvsQ1QffZq3rp+rFqfC7BZooxoEiCqZcGT7T1BgUo4u9rJFG7cxDj1oPRGn8VO
Ibq2a3QSV9sw1w+tq6lw2URQVGBgY+d8lF2+W+58h9IKDgjKy79sN2pCGHhStSWL
buk/w8pv2B3Rotpca2Aodh7vaQK6IMzqH/o2kKQy6uJw5x1VK8UPaUcdqhQJltff
PGMV9sR9v69OXp64he2AJU4ZNwYeyKfE2ni1Hb85hE9Tgs4J3z9H0r+RRthKeAXr
TsMkugszs0zkqiJhBQ6g2rPSKDQZa5vjzkJ5i6KHcwbyGmgV1JyVtXwJh96oXtg/
tj0pZeFChM9RJKwfAa3qnXo5qRIEQ0Jg5RGBT0aWzm4L1uLi1igSpO7biUcuiAO3
oegwmM+EZa39IqmrUlVWQk/Fkjs0HzwBfMbeYgFqxCZCx2lnNRM7oPdIln0NFOUe
+izjtRCUlkYntjv5pnnuRDXWlTANcPIo2pki0ZYgBAYVPfIV0P+2Gtz/D9N6XWLm
kqOXSeS3iNlkYzj97jYcpfIywPIWWnP06wSGL17fX1VRQjbLWYsDJFarhLGf191z
SiGG78W6p7768HGLxS3i9GWyoCBdsBe1DiQoqBKGMXUW4zSzcSnDr5xy6N8VSNwF
ON1H2e8koeihF7MTyhgQnOLh5udftLILjhg6fYfCv+c+OSsPDuQigL59KXKF9AUe
fYgrw4bjaWa8/9zJxiOsgWoYXoUIsB9izWBLcyA1Wdyj322Jzq+cQ5IT4bRJqVkr
iGSC2VhgePvArrDlLiTMtI9952DSjDGzDkhiFrY2X21o1vqAkz4Y0WjoCCoKZ9bF
DhxuuB8Rz3vANKsKb2ODr1kdOo4UFr0AnNgWgdxd9snoEqm90R25rC5YfQ0rk5kH
AwJZ8AfTSzJlvkqvBRzOy9wjmqpikWWC3ZEPIS9VBoBKlgJT6Dn15OL4wg3YkbVF
iRl2yTOmUeVeaxIqKRoxeT0R3EDikfYGI4lNtz2oWS43Wy98tGIYXgMEISwsDyPd
r3J021HWR1xkJ/2gG3iI0iZ80q27xhU88oFVZ+7JYWv7sgDhC5sGK9UG1LItHRES
98+eekc8S/cKdfY4Fz1cFDyWKo74XgiboQGCpIbKaVQgTx2+b9hd0pWItcoYFvJL
btj2c5PLJRrildh+QCoaWFeAo1ASLueO8k2Ume95X+DgG1q3SwYU0PfhIRUOjI0I
HPAttGPs205L3lX6cGFOiidNwK1KDqaXpi0/xTupEcQpSEyfn9jd1CL66o4WiP6/
QflRuq8pOp+JTYzcpLtb3/7x17r4APPBpG3PVWUswD8rrGg/eVDvbv9NTnFQrjPl
cfBH7KnEcR1FPYy6/WaGh75R5tpeFBv7vIPgdxWoaq7bi44LA4ZklnCc9mG742f8
oKNLjoHWN3eTGpsCyBZMz35KWFhah6tIOG8OjAE5HKpqntjWG4ij2+7FO/9PqBHC
D5+j+AqxYcJUHgrkl0rBCHnRxeuLX70QavOqv7s5iKTWM7z5QyDtvJwgJN16OVBn
PewffsRknPBEQW/gnlFQNqMPYhvcDhSC8LqKGM3eVmhhQXe/Fo1l+PkuJYk3Nkrn
RdQUPZckuXZi3njKOggYzkYwZmLo7InFNNgvDxCPsVvuwRSBY3nZ5V4GY/A1SDCI
FDLmZlw5eG3GVS6003mO6lIZXOmBY6+lKVVrm131vRFvi75mYZyRAGWinI76au9Y
ZGGTa8JqpVYXShz6IN5PWje0AF7nxSzqvIIq0TLUdTIKWBESwDpM0I+vGeLFzCr2
fV4tIBnb3kjf8jdHa1jOEo+w8tJVI3239kVJwiu2OEpKP7zkqUS8MfMN+Gq1YGK5
BqTUFcIbqfjOtgDNMblRCzhQ4ASUm2PmIi7aiLeHgYZSB20v28Ugr+zn0hRcclu1
pfIgxsr88/ymhNPZVlzeUTnacI72YvHDJwFDRKdbKsW8PtoSDh6WNGEhyhvJtHS1
6YRzJ66cP64UpQTZQlaSmiHaFgVKzPBQiyCJ5P2zu7jR/SL/+p3sLB8x8z+lQHlv
uozbD8yE4W1vNQqE8q5e3engVjdsyWn1NJaUh8tNkJ81/llqN4bIUmZH61gnC7+z
RQL6rXdyO5tc9MFce+xLt3UBnQvpQI0m2Ffljuzahq1AssWY6R99Y/tsXJCfNN2o
R4ur/P88aEeCXBVedgzeIKZosMovF75bwyTNUmiJi69iDsZ/APdGUyBaTBG3j+fH
yKKSt5ePn+G5nenhtoCUaWPu/XdwF2RgNzh8+sBNlWGdorsCcdIJqjTYXHk3Tkmg
50dWhtiQxv9o0Jud67QJHAQzOsJ18VdJKnO472d++3U5yCtmnFQyQlunTJJoCrAV
AgSyTF7NTK8VtSZb2t851SDuaINnRyM/fy4gmZ16RWP1HQj35d6jpkQjTJt/x/ce
0E1OQ+apXQmDuCaRjzh6HWmTSgTsg3OfM9IaZiMjmmPsP4RLucS9DLQWwbwCg0t+
2AEE1NGxx+EdDsZuskff0UnS6dkO0jrVeXuU5GwbsSuJt6aWra6PdwT71b+oCNfZ
qGxMTP+rBYfBJMjSUZzY/V7J5u5QeE5kbxxQtrT0PbL8FYCm3s4dvemok4/cjM2s
DuTYIEwDMxOpg28AuOSiOX+cWmvokDF/oSVlgc9MSybGFj3vAkyi/sl1FFUF6FSC
DKFdrwjJhaojpUtOGiCmxDRIjduX7IVj/+ANIqpDNkotjqapRY7zwzdoke9iOtIW
ptPmyGjTrKH5sQKqlhuGPar0K5LoL6onSeQi8JdA//uYMMBTL0hwddkXFsf8sd+K
erUCYmZjIPDTNbp06zn63AXkwqScxDuWK9tcteNKHNqH9oXADpmGscJJza1aJNug
xK6rUwZgPEMBbuOFSEvj0bEIpr8k9porNS69VnZBkW7rgh/x2Id1TNK8FdneyQ5q
UbaemDzqMSutbXk7St9mkDL5XwYReTEdBlYz0CV7D5ksLO8LvZkCTsahdRHtPAKp
YBJpKt1Hmr6YU1ZUphIHn2Ppxz59TgQTRvj0d20ZEASPAq1fo7LTbZu8J8RQiVEp
PxNg3wbosaPXsAaYjWgszPuB3ROumKm5cHv3b0PT/pjGyo4iGoDAq9tb7ejevMrz
ntRJV8y0ZtTyWMYKY+jbsSHYgUeZP/6zKL6msxu0naTs4Bq+DSvUSUX77vGg+FtU
Nr7gaEvJcCjLM5PFsiOcyZS0Oqfc9VQWAivyjHlK6N11DoR9UtVnraTUriGkJ/Ug
rF0tasZaIMj98feKbBjfQy9Ybzfn6cekefOTR3Pw1hlZFs2BEIdl4a7e83dtAYcB
APHK3GW7QKmxUHuubB2rPCPH3SxT0SEkBMLQh1e3GGx+XqRPOGKPESmy2ExVwM1t
jbfglyT2w3por78DiCfQAcfEUj3kmVwRJOgfbmF12Lzwf5FGzVjLbF9ka0zCdja4
6DrG6iojlP0R9qTlZEwKztPB1diamQ6RSNEZKhJQ6Uh36g8QIuEXBH27ho8FSal0
3uUlZnlI6LGUOQH+JHTm7CIjoqm+UgcfVRuZ3itWdt+vzbG4GryPhgHKSJ7IhgJ8
+RnGVL8IyezmBxX/THWEIBDXKsu4YaB87QPM+SjPjlIR8N73Fa6HGy0Z8u43s8uX
o93EXRErJK4jxg7FIc8K9F9hhhn5ZEm0pxX8IaGJzG2aoyGKm4wLz28Nu6vPJexh
61WtC2H7+ZIc3PIYPsqAzFpiXKwjbrCE8n7FZyS1JUE2ElirlCZ7lpIknHrN0MdW
XFHT6STSObrJCM9R0KhJ+TGR5+o9I5rC041sWALILoW3+1El6gtIm/LoQ1EHTA8d
w7Q0xfwZ0a74CsWI84jlV5UDg+I8OGenqWmn6pMrpYIRezHH/Gp4jdlkGmVWZsIn
Hf7jkEzYPBzmcT+dX1OdB6jIzDsFId7g8M+/78QAVXj/iKURtMZbnkzpn5bcgPAH
LwORMgpanGzojhQZ9iyywEgBB0uVKS9fJbewSpfarNaU4nEtosGROBPZbeYQBPMT
KBmjaMq3SSsSviGsbcg5DVw4otiQFOfZSECpXTBj5XRwkNlOb2/vWGf7UWMlrhQS
OIorUpNEMPfepjPx+B6+xgHRjM1BKjjMDdAkSFjYf7vtYZsb0N/iXIKFw+JS4AYZ
vjpCTh2Zh7NmS4cJRA02qz85SMGkkH0+qS7hp0mci0dAQ0D768xFnU0ECK3vy/0g
4tlrkBWJNb50mxoKNjM9FbKArBy576zlmtRszLnIZqItPovlvd3guePOSHvqZ5N0
gzubcbb6yV69H+PsnnJsjqVrll0DdL8JGFHG6SwimEBqRc1LwdnDKAcVBde+rPJI
VEnyrVv2DGj+a6I4Mn9rOCukcg25aCJWhx/HbBatvr8V1hHWlH6CiarBRn8yFQdD
QbuH8tAyOjDzFxU7GJWKh+Sckt1EnUK0X2HTgBpx1ITyetyY8E4Up+ADBEQqFlT5
x+QoxQWZRtt5gXptU+Va161EoDNksaQmcW3CEpp0vRhkQkOaaGvDJyfqreH90SVV
SE7CgRmE8go3WiYjQf0T9gzIUrwizNvg26R1DaBiJid/4h4GCtdEfNPrQS1KUgj+
2mk6kZq8HmURMCR/3dmpOmcwcEHlyMgLFVbtXGwA/XMbu57ejeIlwwyUdxCUfKE/
zUbfiRB4rhyr9b0wKFuDC3oTtwHg9labQSqHYGlNK1K6WtUVVJrzsGdOPaVdxYum
VaXILuMGI3L27wBkLLRe8fUZwM8GQiU+MwfXvvktyxntWVc0HZCxwF1ujp8JljiZ
pDJJR6y0jiWxIRK9r0B0nyVSf4+YLoOXYyKCW20KJmBi0a78e38hG/nvybf2riED
DQYbeEsTIYfbr8FOmHPNJJzS9kkT1/DudxPYzbWy/958cJ6HDp3d7izHyp2tgQit
Q8efVC9qX61EvK3khbC5PgRv+RwYfD+3BE525JksEy0D7S5Kd1uVuUXHss/05qDA
u1KE5yn1AhSdVz6k3uaTyHQuLdAQiu6bjR5g9oaBOy6RD4ncu+yn3B4vYQrywiXW
5dnGi+VuYj/zE4GAPZPyEwLQ5WKQDZb5b/DEw2e9dNzfzqlfZwON4K9WSfzk7G5h
F0cYRe8PvhvU098o8OSxn0XJYZNd9DP6ZGW5OQHA2x9u1fEgOu8GuamVn9KZC1Hc
lZ6CN8CTTQ9Jul4zMhK5T3qf5+E2eM0F8SJvObbaKsrnYietnEWZvZ5YH+H2wtlw
6fk53oN6rqSbCE+v0O3EYWBckLA9zuwx8x+XIRtgiCb2pGLLy50fJdWlPoixsrOW
qKHedY6Eozr6Do1yNrsauX6s2+YzG/JWrDp/OCDTnbYEQnbNdR6Mi1tjnOJ7tMx4
We7bDgalkoJFUEhkCpVLd+VHOcp6Em755J6KtVFJWY9IRxHkIu5O++aoJM6gvJGB
UtjbM0z5kswtyJHsm6GJHPC+mW/E0M+PQq8ejZqFJe+JGyo9YIbig8qJvPTebQAb
rakd/c0roMMvTgvaA9b9DX/ESYHmkaJnH46osoFeX8+EHneKpOpMS5pmds252lqY
Y9pAoPebqxD3oFSoSmC0Eo55W5Ntyul/tTqexh23H1dgwG7Cg9B9D38+lrJO6OhR
+nPBd2ulXnrMMYa7ABlTYSd6EUYjYCMnyyW7SnYxoFVra/1LE5xP3n/GUmq7q801
k51+7gZgx0Xkq+k6iF6zYIWnWC9oKb6gvqyJ4XhlE503Lw1O53HoaljuNikNtgjg
xs9YgNmqzpNexzmPS9ztoTj8J4tpe/6u+G2qQv52KMSF8TfE1hX3eUl6XnBZt+T4
0LD/NCm/vuVrn3RfyEjgi9bU4XtKqTxytLM5v5yVbohFfBkk5E+0+ylv95ZtWLlf
NbsyAHAlA+WQKoBANL9rAIhIGndQYNUEZsBuyFzxTJ8KBJdQ7CJV4h+AklWVfLAk
dttdNrvSRyXTAQB4q3uriOy1hQ650O9eqGw1EcY0Gu3uqAFv5y8glQ2xEVZKZ5KL
rQ70hGfEVUvFoSzYYVZFdiN2O3H6WMD4B0xZ3Q/syL1JzfIps/W405RmgsCKfPsK
5gCvDmn2NgoyFkkxE+UP1iWGzTKwVvWnUDXF3Ot/DmGshtQRG3keRCW7hIzJhQOl
7FbdlwoOb+8HiKak3zhZFIutJttdx6A+YhKqi2fRBjq93kBVfsqjSKEyy8a3Lwwd
rZXc89d3cmSY9uq8KIpZwdM1doj9Qy6XE8tCBlV0tc83s5lQZO3tQpFAH7GVc9fu
s2EMZPjOHewyT7grUU6k9iy7iCoijej9UKUSg6Rkwau8VCXLqts5jb8WgJEIlI+o
527qYcYjZrcfbyIexL7yLDSl1/bXq21AzJZqAWIjN8Xr4vg5RAoaEnHzwKnauo6U
xGzVI1WH4B/Wu33WX4dGQ1Dk1pilzn21vwQU/US42MJJYjP/37dA9Wbr3RdHb4om
KA4FmZ+4Mm03WPezE1Ah1tP0Cc6v+IGiMkKwFR5oxQdUrn2nVsDsk3yGeDzyGaX0
WHzF4Kp+vjuPzCeW26EWMO3sGLS4R2PFYBlBhNL30ZbGkHQE/1Q3okPLT1hcUsOb
iNFTkTFCP5gnujF7OVZDr+cv/l0AvdaxbSgU5Oqx0MNePwrFF8CZAkFACw9+CQSp
SL4LYntj3lkEYOe3Z1yEprTEamDBQRs0oiJbVIp5XPu3cYSJ9B8uTtzIqcIoFzKE
NaRfD/L1ZEih+arLXVtwzFlWgDoFFKjneIFbcb40KN/TBBW+pp1Fc+E/VbuXylCD
KLFTV4FQbHrRS8g7840Pj/cHEFqhsNaSZmNTJ78MngR5SB7AXJBUq7ab9hhR/JFA
UC3ONCxDF19RSNhM0InPbXE5D0UVqWrtPgHG2TPY/1ztxRiZy5qwQ9IPQpo8xBBE
efee8Q+/6YT2g9IWn+dC9iS0ek84shOk/5cLjMZQWT/1OMzREB2EKzd3X8GEziHz
jOtZbb1WDsOPZLMDEogXcZRWAzY5vAMW2wBIimljCkaYuvz7F2Xocz6WB2U0Ze40
XQthxaxiJfTMi6ughIXA3bnYvGyfmYQcZjUV/aFprQTwJiPDa9Bc+ebskuNOkIWr
wv+yji4VX2gD92Y7UvpEyspjbzctbkuR8ZcwUet6BXR0A9KICLETTF8/0rvxA5Ve
HM6z0ayfNI65Tfpc6hm/csaDe//5TDP+o52B6Bny8a+OdUsML6/xNT8qw284rDfS
xxJJRY6PutLHCwSZEpI92g/AgqVc1ViqDzFl4I50N7jh478R9b5n1CSEcEQ+mes8
fgl4mCgQOdwKSrp5yyZrFUaQ0K8oYrEp+hfbnNjTW1Op529fK5sF44XxOMCrbRZe
x7rqhwJEjmgBWfN1qT66xwsf6ZkCEv6muP+wZYVamYITjUciWm9mlpnTBONM+tIi
Wh7/NtR8rUssF+VZ2Xnif/p2TM0pBH8i625huzOoJK3jtbeZorKhuthhMu/yJJ2a
THX//8Dl+C3ymHlzMqNMat0aNuiImug7PiTegpl7v9QksWx6q/FyEjTcVv0eLaKY
YqWzZuju4CnFddFqA9YgN4qx4xwf0wDlECKNCF03WhxqAkrA3P4TKU9EOK9pDR9S
IH7zCSatMyGwd+CsEkuWqp8SM02JTzg0vWJOMfXoiOCHY5cqBVzJYUXndVHbkDKG
GSdLKPg/+SfaOOw9UAy4GpKbv8wsx7Fq1aUCFwHNk+ktkS0GZR7xBj2uqzI+QJ7g
6u3amj3KNAtv5LBWKXUiL6qMQbKPL7P41Z2fbLzqtpTvVowPISOaU2mMmQk3o3A3
iSs/XkdrHnOPWpQUw6pt9C14B5Ie5kywn6iQUNm/hZ6py3xIGDJM4VR8/3d6EhmB
u4C1gUkUQXa6rmPbzDcj6+G4v6eqVVU5O4wVtU4lNCe1zETKvEdefo8O9MsaGmY3
SjE/bLP0ebgKlU15N4okDiY8/4aXhgefBQellZbI8sY1DAfUEwrrcVcYkh4wrm+I
059vTwbk+huXXExo6EzKMJuMBZORcMD40bYQ1Af7FGOaZtcoBY6xAlxBKfbh3tv2
O6o+XBhWakD65sYLTV1HZYap3FhBos/rKqex+rVyg7c+wwOHZnE+4Hym1mCDYsSe
OgG4A6Y0OvEgDBWknbapchdFw39gTZoq36ByJzfecRm1aHpZ1RnDoa7E7rx4O1TT
CQOiHOTek2+e0qqIdaWfRuWbh+Ad+vQwvnArYKZdEzPxm6c+ooyZq9NLjaozoIBt
vDa/vmqhndK4NBDY1fjF4rIq5wfmJ9GbKb+ncXJD+8GrQyOi5HXaeDcIpwc4+MRA
qJrZs6x10EcrU8U1whNXd4mjv6UL4XpBx2Xz+xCJO15ydjTcEs3jxezeGb3rEG6f
6SBCMGJYA4gBvM+Eb2xDEecQ+H0661WXY8U/zTL/nJXy0QaSB4z5mz0vBeRwhhE8
YePP77liFX3J2mLRZT2tDL09JC1r8FAkQgR/qrow9PT5UKl+jBhuy5BciDqp07gT
63/XoxAwwvnX32cq6CjnQ9bNvyfqHPITZ86HJK+uvfAUIQKCvbFI1XUOulsRiNzL
ldbQoSGyViEThQEQRXPiDtzR9rBXbSYCkcjwI8MlTkAs4C/uePR7MwfhhbjCGF91
xSij1GW62J21akwz9kp3sJpgZlqEhZlxGQIERBE4bN6nwXyKqlVtcN+R3g3y5Cax
/tiBKgKcmn4NuPKrK2I2wmUXiUPR2eKZytaJulpialSaLyYLvvB/vdk9QN6Mks2g
rOSB+lt+CnOqMaeybfpJVNAmgk2Q60TqPe/uiYhk3L3lCauq0LMWYecq5jB7IfOF
jIpuW8+orlDLS6zcgxlKQe6bf/Mql1jiA/GWJgyEDDdRkQYzBZaVC3BCtMQ9iqSs
H1B8MGL8p1/DWc+0k0HxeWHC13c73XZuBx5yLYyFqdaBP0fDOCskmuEiYmP6uQ6U
/igB8fBIp2id4NB2HGoQiLyCoFF1tkAba8O60neTyVWGwx/iLSG1TVCj9Z9oZkc3
SdhM3bkKwRrexqzABH1IFUvQkYXRF+GdAqhJvlLsg2WqUeLHk/ZNrnqhfJSYUaVO
OLznNrllh4m6UhzFJ//9zeYGml1rXOfpLcBbRIcVXWeur2r2KC1AsbVEAzWqX9mc
B/yVrbu06D+hz/kgcQUADgMpECCz294Lg1i5g6q3cQcJcIniyT2CLxMbqA21BMTD
mFCEYN0bxVQ0m3/mso5meNrnn2+iDoXzhzqo60P+EtQqrZee9bFo+bSvjeHODQO6
QrtggjR0BBwHrGkOLjoLa5hZ0nzKfWiGtMlUtCcrEWy8sol2B/3emHMxs0ilUJim
fhzFt9G2DJ3pTYq84mjrqN31smnBXThs2A9xadO59h35xmZ6Kqtj2qrWTpg7kwFe
TEZmhzxZige23jwAWwbZ+FZX/mUcl+8+0NoS0cman+0fcUrINKwHRrGUJQQu+L1c
Y7+0jsK2q+r89+a1VqKIP5+KOWtJ3tbZunX+x9Q/vqVOKlrpyrjYaUueVzotJJyv
lQIihw6MLwNvtStPd/k/O0T5dKqcKfNQgkTE1MqvO+P+6nYOrifoBOR/p/C/UvIV
9Sb7PfPAWyXVPsxlcG5jyJnBiMlnHzep96Qu5jEjQDCsGG6b+oAA1Q+tXyTylGo7
TLJ+7UXBHOpqiYSdEVgArFnjzV452pmSUI3D8ojK0oh2164TENQD9bB/dMScfm7B
gd/cNMU5B8v5B1Lbxf4bdDARr4Te0eor08hPokR7PyVdbA0BBT0vaouyfad5tGat
0KdtFQd/0feg5/g00TQb8qq2lp3Le7suYdQU3Au08g+belHTdAAf9B1HnUCMAm2t
hme6K1yOrvQOZzfufUzvQHjSaSweHwbmIKGwIYYuFu3kPr5VufoU5cCmS5kKPVo7
TgKjmdM8k7HkGolcdsuE2Wejf+356ahBWTLJjUurTncTGufLp8BCMWGhMroAvwZM
PBViqnD5JUL1p8cU+A6odS2rH8pTZ5Nc2CKpcoG6YHZ1+o9KGFobhh0awtNb5FSY
J8ROIzB1UtB5E7cisCb/IAu373EiDteqsVcuk8+KC8LnA1A9jKxGYhLktADOhOR0
atmXrdvCVkksSQhR6y/gxBc7hLEydmU+wKKowdVb5D8jU9rR98BdPw0xGt8zmfU3
5uplTFmJU4sUkDqgdU9YEE93WMvtK8gh3/qWihd2nXGn+sUbQ54MBSFS73SDHXJL
YRcf1RPaRSwiPQb4DR6BnE7kSxGRlKO/8NUzI56Aj4ttDEdoEmLIg3IP28FZNPYS
qNCX+5qSVssxmIrlgCy4KzwHIDcBpUR6jLaxPPIjKtlnhLYKKnHAbSDoBN0cYwJu
LRNwss/nyVpSR/CgWFh1a09VSK8Oeb1qSHjjGZDtgrV9rTcyRPf6MvASDHe1st9+
DsSY5yIbzOAP68XDaW814khoKFM5mBUYxQ71QybhUgJfLGtDee+fsSgOsd18meXu
SRrTRbH4JYmA2h4WlqCUAPcHERP9wvz0kFxs6i5l0qdPh71u+hrS8Eca41MonqPB
zho7GrrQ/6N1oz7Ac1HCPryHL6kFFiwg5VI6yzds4wJS8FBAubjQpVum6JWsLdln
PO7M/5/HcfPCm51KioNpFHb5R3ibfx33Mg70KSA23b34zQ+dEl9IM3PM31RegPSS
YjVPpnE571Nhmz50qhXEusxZuJm1AHxuh1iMmyMieO1gMUYRwJCI6vvm+uuOPEfq
gtYqnjSMvPaayaMXfRxvtHrNX8pb9pXGFhWCofWfyWUkkB2mhtY3BvckN6bUWHK1
VAIqWGaUCvPLCYIAo5Vb4Ns2wgxvhoTFWx4Na7u/EUjC+WIa0sIGEdJNVVtBgpzf
vWVlROarIt0NqZqctR95ofSFihl7eCXmexkwgRoKRvbeJg2Y4BdtzmJnp2CHvkPj
6CJpNCGYU5jRixCjmNDfEBb9gUBFaijzElDVsvc9XGZawNuS6viBcwTd4AbUqsQP
qGZ+wbSPaz8QPxmaC69/Tv5qncUyRBLQOGdpl/+nM0v+F96dIfPed3BNaZqMyk0B
WstTZIydex/Ee5Tv470coQoz63haViacNJ9QGutCI5WKrkZ5vhG+sTJ3AzOEqcM7
sNl7/031V59vIjXhhtzbukLO6byS/Yts+M/JhZgsu5MftvnOqFcggJrd+IIJsy25
heS3rOMp1PBSMxR1p6UEV/yO/75cRdFnZDq1Ke1ArUAxWfXK+Hdfwy423U2l0MNN
jVIUvmiCjUZrlJdBpVKs3UTBaK0mZbo7xQNCaW05w3HL3kBo7020yConLv2xopE1
OKoVgJbHX9sUZk0sGRFg5TyPPMZx0PLZ3/DGX22UXwXY37Peg9bFAK5wFXvm+FHw
cIY0QYK5bWGEnlPEdY1eGqzrj5D3V+Yn78gERDexO1ndFy3uSlxhMv1NfOoU8vnO
gbqfU3OAUPMcRfm/Fc4TwKDHYrMGPKpLuvCzEeSAOTmVUHhxO6c5HqRDpjD682Ts
QkJkMuhcOB1MJn+QSnH7F5bRE29w8fhghs4jTiRiw55qzwYTpVLwx2KO5A+YFEwW
RBnidjNxhm9xsEyGJ132GGo5VTeZHt/86RNBWDnRi6GHqmG1+aA4lVSrVyThg/Fq
FCjBCYiJhLjZ/o8fRl/KD2VMWKTZyK7eK5ZCtuJR7xb6Q2AZrc//+kh59K4eys4T
3nwme6NLIt0lbVlPlmhpFCtwwpSZzfwszR1lOSoSeKyQXjiFz2bfO4vR/FpvKc3I
buAgMjBpUX/7W2xZx8xUgbyiEK6Nm2EG5j+ckUN9r5OF2KdoNT/wHsPQbwIeEThH
ad+K9gEBhSl6D63EwWnQOL31pzfJgCrl/iuDkAeORLE0NEtlPEY0FgKSWYqavTzi
R1Ki/2Vr7uscGrcG0piNbyCLDNji5PRlvRUrlDclHGMpwLY6HytTQ64RwCKUzDw9
9iSAJKZepwIN5nR7518mimsImobrILchLq3HUNNhj37MlA96b1rl+IVmK0RbLoic
R2OQSQv67lt2w8rJbSPj36LoSNQNUeoLpWreNEhI9WKR2EOr6Wk5JRJHm8P1ekuK
cR9ds116uJM9WltzScz3pWQtHNAHvkZDJz18fVFlgUCEWzKNbsh2YOCTmNGFWYJF
UM1DEx0gD7bd2ayXrQa/Vss6/72Hu1Q50PXXOo9C1x2ArIVIlPxT9BRm38D62loC
uOSJTk8d6RbGkzIIq/IR0+qeyZoh1POPgHjm58tyI5ygATD5N7HC397OS2kqAIVo
Iz/6uRj3qDJqMSDicTdQQsy+jorfxSmWjChxSHmFmSI4zVTzvmv7sIJ6nQGsgtq/
bqF4NE3MUF/FOL5+7jgvM1l1Rufd3DqHiLRjceV8nVs7oWjCHkIq+tp7qVEVYvNh
JOePi3E/hi2WdIef1WEspsQzX+5o72Q626fR0sL5TRgaoU2Qcp/R5zWsOYnsnG00
w9GQ7hldMjv0mBi6s8VSR/SgFL6C0AMJeqP42kzlVGZAhzXVycBLkH9m47o+/3Qx
OXfRxWwW32RJoa2dnnElZ28zEsAoO2j/bABGTFDjX2HXMV/7wI67x1JN9TgEMp/Y
7PSQkNUQ7SyMyu9Ev4e0rmn0VvC4JG7ds1u1B4tM2l83g0IHOf+Y++NeRWql89UO
UNJ6hd55LHACChp8PdhAxr25kiSPFQJuAAEdT9tWF0twKLok9U64g7jha0KER7nk
DGQCMw2c4uTPz2ykgb0SIOihw+qiv+Aeg22C5wVC9fEa4tX65qbYa9T6LkfGXiRO
LY8zGBhfgmldv1D1Ue7YupR7Gq3WWmCuEZIKDLGeXQ17kL52A6jpImJdJkxmXC6n
wrE9uuJtpr/QmU1VUU/cGxgnAKxT6E//wf4+9Ew43pqLeHwool2cxsx38y7BXn7r
sLz0FK5D7SD+3kTckfCPmpOaYuplesH4CGO+tqk6/J9s2yuwzUxEvMydzYhRMNYI
QaI9M0PqxxkKpLrHu41apxypOsLvC9S/1TqcjEl+WD3/1osU6Uw6yMiFXsfmY/Zy
7FWOO6AF6Xg21yIpcjAVwpks3IWm5edBDsMimndtvF/OUTDhSYmU+XhRN+0Gqvr3
orlDsyWPVU9dHvilXAxR4ydH+dhb3P/5L/UKyFwQFj68GOrSF9DDGsR4vwsGt8SN
h2d0Rk+YFfSDzpYeicU4cOZoxnD2MSaPK5AUFOPMwqqYTtOxPB4gLxRC9gLiLZs7
0Zq4ttK1YvaiQJJ8H3Xrh9XFDJmCAvwDCvssU9prISeaA3t8mznHWnMqAF/0LvIb
zbA+RRmLcHiyfsVjSTiGU38d0PEc4idV8G9SWUhRWHfv0GLD1KFueU8M60qRVcVw
WHesHMA2tHqSCuRJmX2+Nda2xNBMhL4Z0oa00bO14bq2oDYz9dWWwm+lp1cZ8zk2
O6flWZPS9ozHfZNRR3WxnMvsaIDHQ0lXn5h/IQFMUJxa1aGS6BEuRUD6Rh9iKt2f
ZOHd/v3mm96hSMph1Sl/2wFd7SKylv7ywn9BMNzcNjccsO+xhvOxlrQiraeSVGF8
P7LwZDMhe7uRMRzh139YeIjaU6Sd06QAqm7IBqYyU6MSGiouX5BmtQeVkAx2r4Sb
wVfitAdhsSdBZM18r7uQkSt7zmSJ1ieRYdS8vPOj/yp+vNdCpxL3FZpnzsd9JF3c
pGDpjSU70vyOy+m4kqLs1L5sQQ0Dq9HyG88gJChXilNdNJHYEAmGUXDOWbQO7+a6
sQsK7TyKJy3gKt138ja63GOzhGFEhCupONcpJbIhFEMfiy5iC46kQwL6JhM1vcv3
eeMeJQvsID1Dp/DuZWQFuElBUSvv0uEtuQrphZrYhoUu2FCXhqKsPoirodY1hCMv
UnaOzRMDap9gpBDjnJNywjCiJYsE2LuVYoqJWGLSm0nrErRPJBQTnGSRNuM7SO99
MkmASFGBRCIn5uk2kNHnPccwNh30Dy5fwzNQHJzSe6k0lpJxw99BCXS4v9g9QsYL
nrDrbgVGQhEMv5RdT5fzWgfurCRGpfrptgvMKmiISBCXOv2+yJmLuC9Rgg+NTTsx
FX0pvrV8OA9K8tpCfmycPz5mcU/Abs/yoq2ukbI0R5NNEylRBbQC0jaZ++/Xr8oe
0Et3Di7DqirVLzUC1Eqj/JDD1fBBQonHuw7vExQtkiYKYbs13DjkFhyJoc9Q7GXe
M6x9uecVELdEiysazAw/pWe61QVu+Sdv+HkcjTXQWAZ8ZIbJkCNY8UtNRjpHcc67
2VjtQeH8hB0ZYTKCu5Fst/tazHZ7gav90Xmk6BnA6Kb3eEwd8Hiih9YVMsnHyjSD
kEYkdv1KLdFnPRKxhEwXxniGJHLoJBq/dZPt7Fo46egz7JnNqPe0brZ1iloFlXHC
K/ms2K+PZAk+FtDJb/vfZydqoWsH8AzJriO35vAP4VCxGnMWTlMYBqpnPTLdRCt7
G5kVexLZMh7rXF7JXCqZXhzZ38luIcf2kj6U8WYgCh/5ygPJ9z/flDblMXEF+PPR
86vmcTnzGsMe/s6jT6GMMCyBwBXJID7phM6W+4TIZ3C/Sx4/ERoXTaA9wbbe2J7e
KeuPjYqvvumNNx+hu58PlzcgOO3XgmKLHIov+cY1fSYYaFARpsVQpVKyShAeGppv
uYy6vJmGynNWJ3Wr6SNLqKmHsY6NErQUAkeyo/n7BBB1IbN1KKaHbuLQUdrFeSYD
lIL3NQ8DbORzbmMzNUADtwjGVcslOrv+rzwz4LKsDRSs6C1dgoXPeZFM2ShCzkIq
e8Xq7i+3/afwQxsPTFtkKR7rXprZeU+WbOmdSCfzyIun5CnAiIHsUNJ1L97Ykvq0
5dnHGjg4iCH2gJ75p1UdeLLLxb9y95TsxTM2M/qxvEShGTOcInd77Z56Gkrab0/l
MYpoEz1OqusKKfP8b4Sap+eNAQA/wUNCQ6GExSITR2o/qyHVTCp9IpptpV6/rNi3
h8G6/9gZ650ng8ETjmvKIt7+saI7djWQvyjlaQF61f5ivAy/cJFJlUfVmdggKC1F
bTVyYguRDFEOftTkBiytS1m3+Bn8anz58akNzckmrLIK+vTC96qB4q+FPZ5xAtNJ
syxGxryorLhw+5cGIR5OtT/jJs8rZk7WKuZkYrUaOx+++jT6e3jJSJamAZNq/Bww
Jh3g1PbQ4bwhqVYGmiSChSilr4r+kOg0SNM76rQhmbbOcVLlPa8zP5B41PYtGBDp
FuATL5agGHqg+HcMpI+GZK9dGpPoMik3n9RbrghN2T1P0AZ30DXeCqyenIWTDMAf
pAemzjZppFF8FSXrVj4sJIbd6guU9lGyOG0hGmhdGN1NrxJC/ga0dz4UiXhiEu1X
lnpGWSvCS7F347E+Lj8axBUbBf7fnGMCY/FFAm/CcBTYr7p1yMx8iQuYXmsW2aK3
c/ADkYWhwy19Te1KoKVuTEvETjZy04MrcRqZj5qPvJ8J7WWVAoWY1o+IlC1c8PNK
/YvZu1ZABvbsvT86GnyVSQ8xqY25z1xbNiobcBAtcX69PRTldSfjK+P2BLe0vJvj
3rIKS1tRRxNxzLwM8hNyul3LG6EQrxZRh0O2RZED8CqzcUsDVSbtCx4Lq0aJzEje
9UDCG8pFcNvqLEAJ+7AC8HwTd6cKkpnHThBUR8+rrHa0fXHrZpixCpE3o244c4pv
qTGX5xrsz7YniZUv8iaTLUIYavncYreQkbiR4zfy31aaJHWw+Nojnb6L/wqLuRdw
bWuZxZZdb0aKjLAZRFWonScAJ28lcPzvw1IZbZvtJeoRJGf/IRLaIkF8wBDvbsJ4
vr3NVRMoz/fmssaW8yq0JXPuca6dmg01eorymWR64RQB29x0SGRuTPeokonujt3T
GEHecrc4kF9gEhfnanmr2jLTEJCsWwQM5oRUsRSrFthqWCHz0iV0M+oloiW8OfgJ
VgEMVZov+3KM3k7REfNVBt2JraoeeGC8PIJobJmgwo/HZaAgGvdk8gjaU3NomZeB
y2PtcI8jiMhfqhrBpj6uhfy3mWYCZPOrfWpWufFmw4wMqMQbS6GIoLLkHOb0n7vX
dfJ0X4ve5pXklYrLtkHVKjpc42RnyEny4Y7mqg1zPnH1sr9T56AA4OBdf5kPzskv
ejQhxHK8pUHaP1lRIXJGqc2ejlg2Fq/reKqjTXcEw6tMwE3/DeBl1NYt4C9h909x
/J8VJTb1+wGYwwstPtiAJ1+THuYU9dmllBRdeo1rXfVjk9xXZ18p9mAEcXvG9g+6
soPnwWjmynlf/fpVJeu/cWjl7P0lbYnq2pNSX3uJNOqVhyG7g6paC4lCc447G/vU
IPnvNphyaTkvpJ2d5O+gLZtTjTBi87tb8DM6P2aPWt52r4a+17+4A5RMnVz9ny5J
9n3r8eeLv8X4lY9h81jrtzTB0wzV5d3Mp03R2xfeID5Vc7nM4QCUslCxvtkyIW7E
VKUcAdfFedSggfzx4wXkp1SFmXQQMrAwO+c185sdDKSYlMS4ZdDcKCSvgHczmsNu
RvNHdRXUviXT9DgNweWJ6SzH+4NrM8XDZ6BWu1ejYqaxbCt7lsFgMzZR4OCcMKfo
ABNZxxEeqd+Wkhl7Bct+NCDVzdGS3gHYc3T5XYq2NR64pn1e6j6VSajdmYOQSypF
O5nxfA4Mph37Ls6wTxORJ0/SkgGge6KWMd/TZAlEocUrjcRXWxE1Jg6mZ8WialHu
nW0v0zYyrMEJY1vz3bZvzNzm1VzM9F3uTqI0tiv2Q8n0rLOAEjmJCaiz1seqVoMf
+cg4Nd6rnMhl6SHNg5h2zRCAlTa6rLMPAzNSzon/WbFCnHr8ADv1A9rf9baYOGvI
fwEDHdaSCF56HppIZJd3cjYo3NN0g9DLv1mGc5Gu6qsgMh0D8yOW+BCVq8DgiirV
l7S3WVSx3OjqeZycjWRxlGEaY+Sy8vkhNJj+gEMT40lupGI3WY/r89STfzxyahFb
3++RkagJH3dYaRxlgDYA53tu/7bSuAFXSEm3UW/RycXmtNTmO99Dd0aaH4duIWKb
btHiQ+IdWswNeHDY293rjPlWOPDzPpaoPR0XJUlQE8u6Ih49eY3kIqCPmipFbhib
Lrlq/HongT0OMxqcSzpEk98HULFzO0eBV8jLXf/hVMf23SIYT+WEx969br17w+5+
Dzm+YWiOAV4wyXNhSAkn31wz3XAfJksNCxkiUt3phJU5oAxUIEkNz0qJso3XKYuB
pGy763kIbulA5TBNTErGPYzrgWMRga9BNjIkC+HgSKvHX9q2ZyPE9juHWbE61BfF
1eFSdD0Yh2wSXIt4X/OlC18YepoUYUuaGDZZZynQgK8OySqiGUBzyvADkP+fhN6p
ZgiOxWAVCPhCca9GHIZj4xGArrpl43LmULAJv1ZAN7hRQku6StS3Ts4TCQeBYhex
uM65SnybWpixkdvga8x9JV3VF04Tl7VNkSNKyWKkesxexAtibuRuSdJhJfLQCtmg
TbWEXRs7ZcwZdgmJbw/BM/ZgUB1WWQPaaspzL5eef2ziWzN7LOjuYKelMiWySVWd
TV6UKjVN8QqdDffif8edAydhOr4hxnopcyQy0kARZufxKvkZD11kav7maxDImvP+
wHeZ9fXVephjhdWAMGOXxPCMgRCP5F1TnrpP333uKuI+2A0ANHRgRP4eP3UKRwS2
voe2e15tze2bp8jdmfoMdNqukK2Ffq9i0jkGJUt/F5uTY0mKolgTZIzOtjdzMYpQ
YgCTTAEYwik11oDfO3RFYD4yvkfqVdRibiEjII8Ww/olvMxfqkwb7pR8apZ/z3CF
SxwWVHScIigfGkMhzUVDYB9gbY8JbbDEOJhuYDHBpsEnS5vmpRslg5Ocfl0MIoiq
Ejt5C0cE7QeBq5R8U2yKP4ukpaS9eMRZQnjD+u2wLBZywNoGQsicQuatWm9+2mqv
Phk5waLgeZFbZGA/542Ci1FHSPuZCbQMedb0IitwhAYuVPHRqvBNTN4lp/RCKyQx
EyzL3Dav0MHNyiQ3LO+jlgpMmj7myHI47ajyubVnqNU61WlzsksK4KU7qp57Vj2P
Nhi4r7rZzcxz5WslZ8DT64n9fWmRcafPfUE5OIZFk1AyQdnO8wHsfco7NFhY9+p9
8ISPNp3/HQHVtcsbX32GLDsJZNwf4pWcvuSJBW22wI2Hzd2dXBEqt9UP6QeFSRP4
asc0IAlKIE+1mJkaRoTHpGCCNl09cr9hzZuBiGVk7Ww+8uIcGQbiryCVw9leNDLM
b6z34lLmNsPHPuls/G1pT6pZXxfjSwppXCnVY5PIdlvZcRHFW2Vl5E01vrYv/0Dh
LlvrkJJreivJsDXpQn7W9vJkpiRU0dZfS96MzKNud5zZmHfhOHBHyYlJ8KxSCg8n
AqueAf5KmvxABET/ooCs6bz93opTjwV6o2eEN0NuC43nK6/K6TCGOnL9Qey+K1Qo
hUqsaoe0pCvVWctwZ6ImH+PijaWITu9HHOvTDASbhwi6GQH57nS56uXrhlK9aTlg
LKnE45Pnnh3R+5okBm8wGvIgEkJ5PEyvTWVMvORSWkTm3S2dLSiVOAfr2AmaZArw
pxmgGATmg1Rypf1o0pofi/Gf+FYwU3dSVEcclgW59qwHF46jXfd+BTHkjGcbMB9R
8OKG9VRyj2T87qCmzrVOJ6y9MWp5dC6Qg2qTTnT83ADT9FIf0i/fN9wrbR7pNlgK
18u6x7UQaTYotYlW+mbwy/DXSw3qB8LgiL8ZCiYtslIy18XxdARj+YMMfrL1/Pah
XRwBrugJK0HNm+t69PuNcH5hl4/vfSJN7c5tdukTMl5tlIegfURjNx+VnzqK2NdK
HCXkQD8NBJLVTn3/4SD7gUYQb81h+y6XFyObCOOEzKmKfP0uhD8zvoBnvh/DdFgx
wlLvCHMoVCGld1kSx7F5I1RnjkkvWFG1kZYmOHhGe7PbdcfqcyM2lTGXfekM+abG
y/v6WjVo9aax0mYwOzcERFdgtP/qVJKFr2dh6q0zWoWv9PHqvudckhOhJPwliQ9M
YM2JURjcX1eE8M2taSDKCTIuiRwPIpCJCLBACe+YqP0UCzbt07l9ooM6IOvgt0Ac
pQmyzUsP1N32JCM+0HDqPW1SRJ51Ch6Tq6uYTEUpz1Y+/AQ4YBkH4/0ntpZ2l3X6
S6ZrKSc3GSNg/s4r5DJeiW4hK5JgH3QbMBQf8jpz99eIt6x8pcl4KwROkkk3Tw4n
aRpWpTTJCG+oyGJfFESqWtqlOdcAzNC8QTobbRP112sAQZKlCwqdl1UoMFSjmBzW
qodCAx1k+49efPEoY8uJNrhV4V+2ZjrW6XCRDhZsgoB+doyPasf/F2Lq1ZUv9n9x
Mg9SBj0HXtPoTuzSI8QHLLcMkHiZc3o6qVqooslRcFvqu/cDjXr3O3lI3A2VAchB
p/kDog4FANtZcfdzzrcv7AUGwyDNdFoqzsJ1/Q9EYBLnrqlZnlWbtnj8dDBArCq3
hOaoSGNjJm7f+3ZcvKRboDWMHhuhLNRJEQh+qTmDq2/47yddFymw9hnZUPupLRWa
sVw9h7FwjpNEVZ5kyDgeSBelMuJS8q450ioAfZ8d3IdvDi2RiW7Zb0eqpp90Rzx/
YzHrZf4WeP9VnGwSnjsNy5yXE+q/TqfXHeF6dnOj8YuWyVRQATjW5xp63h/XCTU+
J582lBctzUQL0aSJLZtTFOK7xVq7RW3ZkZmDmH0XcRz/cdQJgdldd64HW13AIGAK
AhC1Iy3K+O6BC9VqsT56H9R4jFNaCnv28KK/mWx6NmyqeHHFi4m2Jgux3ZRZSAWI
XWZwD7dj8kegr1ehEZyxeWLrL/uSAY2iu/HFuXojqRHSLZoMIjUsmWLfPVbD15YW
swR807Ravsb0r6WB2EATpuvsARGnGoTaCX8nWD4FObXIVD6ahGXHTVzbRsErpRrb
kFGnKRByfoF4Wm1NVzzXKuIyAghPFL1W4n1xJT6iZlpR7UoTbaOMAzjCz8ImlOEd
DiS16GzZLCnwuvHcX5/RyYadaCujDUzoi6t7pC699CM+60r1USyicM4L1v6qzlMq
y2S3lM+fgPdc1BhG2hOx0HfPRmKDBxHRWRGsbwZ0rKD4IYPhygKJ18l3fZz/ySQ0
U8rALexmbProtCNoJyCYYBfmLr+FZBXLShTigK/VLoayQF/1N79TEWA0y22x4CYJ
3pM2lmYD87RMK0rIc1k18iEt5Ac00BYD6rK6S15qhfxIFjwJeCc+1teeW5YZc2vN
6ovDxQtaV1peWYKAFZ0Pjf77FTxhgsfgIBZH+ugBqgA2ZO13eDNJ/sb2Gx+epyap
3ckaBse+gKb4YF+ZJhGMb32LRLk1rcL9GWAUv6bMx5jihDtaiPdRFC5dw4VrqqDp
MPgjCUpKBg5FkrK/OuipBBm0mIYHKmbfE2bBoOAI58dkjbApvQXReNSzltx7UDcF
pnyd20cKdIT33tZ3+Jb8ojBJx1X2MXabEjZ1+PIpSI6Q+D0yyRgsX/MNTPgvCtPA
lGx98X9xp8nkGTzjCUVWRru1Ug8A+ZnklzYRuGgFXk8R08wgUJdTN14bJbo+ipud
VyB95QNUKOM2SFW+QJEe/8vRNxOzAMrmSkqc3EZB9rAo9CVkWCaEawaWu5UVriSQ
pcKCm9qOKOrRFUNF6bUY+Xc3Qcs9+LT4+wlHOf23+yDJgT5JrCNzgQNBn4cAJLlj
zwk/O5dRG5UKwSUoCJcAHWb5Tpm+9NE3nQ2/sNjALMjs1LmrJJEIJax+JqlQ9/q3
ttVxAV/RdGIqT98H6m1EGXLAE4t1YwBvcdwyRsk6WD122qcewnDGl9WRRMyLZ5Qb
q5Keuy6EYDbSlPqWT94oHlYN7uGSS8Idqp8SePNyGRvwsQcZm1gjsQ3FOp2MXIbQ
8TM7Bvfmn6Re/pcsP36ay2EnnkV+v7SoqiEqFBSe6ebGQXbLVDwHTn2WRwbH5oW+
jtZvdI/UjHc3X3CNWL5T4h2pgMbe7tRg0cwFRoqawfZgzMHKGisQeKU0YBTPR5Ef
pwnprOVuEvKBQ0x8d1Dn54Wpw/HMChKmzN7TuQr7sGyA1qmTjfsE2Y+cXmSLd8pr
p4irhjeiqe9YSBhWhg3zqkCvUFwNYN+jKQbHvVK/WzMz/fUQMLaq8AC1GLzm3ZNH
jsR0S0cfkVZWWUNf2RhN48rgJ+N+eDA3J4yRr+00s+mZK65n3U8D0hV8J8udanSW
HWhHV2bIsajbBFspAsMmJgqCS/dT5toN4e6VN7XpQWz0bGGkLqGa3cbZbSPJNRJL
/ZKG4vb7X2itJxJ1EH40XvL3I6OSuxGdifCyfhqoS5c5WKJ/9sya95AB8sOaiS20
EzjJrNzxu/TZKAU5AN/+ORvxaRShifrO6ojP3Q0bY+HooeCX8RVKiyZ2lkaOV9A8
y+LK8kCpjO+us03uYGNO5fNsWJhodzJEA310KWjBo3IWMG78hGBDa8MzBdC9FgDs
p63pbB/sT2CfGxOo09Moy0/I0Q89hEjEvUV9JLzasTXWIFzhSg9M+j/eqo2hvD/q
ijmFgSmWKtRM3TfRkOugvLsFY54eGvHI37yDAO8stIiem7K6oSCn2rVC6UNieU1o
vUchFpfiQgq8WwOZlfGd2tP/+hzcd5HbXrUT5XHb79DnovUlvH18q9jxOS7fzK9y
k1pZLPDkAiXVEW+rqxcMhfxl6bFwJ9Q4F+NqrEnVUEw4VrUfHy/cuDwEs17+nwNo
H+2KI5hY18r5tMVg0I90L1JEXnciqj4mVxZGbqd9zFpBdT3gujN5E+zSzuZ3VfRP
YAzQx5QTAP6ib713anovuDCqgjg6+p5Hd9pHHkmpbkXm7h5fKCiUv6AXerG9YTlM
FzCdsOu7wuVExRLUjo1okXfbN5kNrXgcTMkwmcujy1Hc6WjXTyENwntWIVA2IPim
EK2HBgXIkfWMKqHCnWXSMEwU7+p/oSQIjncBYFetgNwToVLVfLYwV0ltbZInxtFb
oGfv7DnVVjnwe6/qItL5jvw5GAS4hSxOLMogjnr9XcM0u6gYRH+Pw/94t5oyWylr
cwGS2IQ+yNIWYA1WSr0vbzls7oUZyhIqOBhk+xIpIgJmQ1a2zIw6aMPYt8+WymQT
/gt+beloa0JiCDe7DFjF1TgDQGkNPAwiy/WfZ3K4A91DViVsJ9kImbMGkyFj3OnL
vQZBjISlg04KQmyFpL4WJxhgZ4ZixHjUD0fx6kw2dAhRrPpSpbX5GTNYeT/V/Fok
4i4dMmzWP7fTagdKW4Hd+J6BAc8gVl/YhxcIWTNu3epnKrr1WNaiZFpZDsa2AzZ7
uAhBlEtGq2ErM1i7+CSGH5JO3r6E3yijsq6wI40qbWQEOr6/TUGXGnpW5Fv46c/c
iAo+vbjwLImX/O5YjPUiABXxXYFZme5Ue9Pxf8UmLVjL8W1ovJp51772aH9Ff6hP
9HwJChI+eThCLkZMqJP5rAhRQtPcO2NcoLgj38gLcir+9/sSYninhBc2Zi729Jtt
MdJIrAK5ui6tZko5zXMjxYcMOzMvEmR/ndFv06FtAixAJj/IXAtrK5tqp9OMnK43
jlD7ptpeZz64ZohpiBw7Isnp4V6IHmTbiNF/eDDH/knJ2kA6sWIIX8HXsBisTZsZ
HLkexT4Yd8XyqZFjZsVSBkG0T/ktzJG2GutLaXXceVp1BhH2NbWyEjgVxG8m5gGy
00B6dr92f9ds5Kj5UBu7CKFDu7QE8annKSiIXy0AS4HTXK8xzhrcD0XC2yLAQyl9
8kh60YHxOk8e2Iz4s3TboLPjrQQU6bn4BPzpH9cXeYmDHQOp1CwJBnKC43RmsPpC
OhbzrdgEJSi6smVBBsyaltFtOcN82YHyyOLmXBgiOik/xQQaisNZO1tLApnwA3pT
4G1jiJhIw9Mb7KzOim//PpevN31Py/d0UGXzGiGcnWOfQaAXzuus429afSxS+fuy
yTXDMVrRk4vwN3+G/Ai0gB0WzKw+S+AMKBERYLNIPeFxkeT6so+5zrz/iYhgg7v+
KGOA1yjjeiYFqpdbaWGnXgs+GvUy5++ZoNTkAObpFc52M2B/QvOI4Xp6qEYPALSM
XTsPsV8nhK2qmqAK5KC4wgXKvX+V3qCtyIg64LFWXKqEkXQXe2Tmw8k4HEtP+8lg
MyyZ4RPoEq5FkRwCafl3fvIZK7wIDNC2wSs2ib75E+MDFm8AGi7US2sSIwru4QCz
0ay4J096QVTbqWZKQnloLCCfDJ1lG9LPeX0/8RdGuhg2R+DgQMYz9RHfz9n0PdJj
zkOnSS8q3zz2kml5eziOwliCE4eOAB+0HxiBhw2aNIOFOWV4/S19b5KSerxnHxrc
ZHhdcZokRp12l5vQyXxa1Q2gNQHmY0Dlj+Vz3USRTP4oLFJmshXeFw9cj+9eBg9s
l1fDI7rhXVsbGZiX772M9WV6CO2NgA8sCaAdSsY5WkdNvARKdNNXpRFIbwSM+I30
n6bIfeG/1G2uWI1pFQjrYTYVquTixjmljucOc9TknVjipbn4o4NaEIyXWgZtFmt9
nf68IWk91mKfEAO6RO4UaGYRPAfL20JeL3PjU3FL9yUjBsyRQXBkQtD4gQMXWxAo
VklS9O7nsLCAPIMk/9vYRa07HcUJ+CKJT7nlKrl5qe92KihpAgOlxUe5xlIPJEMx
YArMIWhpiKZW/p6sWt9mWN5aeSnhzx6ftQ5Vswa1usNd4gWnv1SzS6nO4V6yGShD
g9/Bug6lMOyq+RXkijZntAc3GrbKbzGuJ/RpV4pozc6FTW58Szhg5OItzTAnz/Sj
4DcnHP5opALEpzLRysD9VBqzxoE/C4Zir9HA1ap5XJ5SG0S03KQvR4plPUfZ79OF
zj0cUPFU6SKsSfzarvJo2y5AXZAIsnHVLEKTAjFuLwLyrBd6n4cLnLXN4yQdT3vI
+UAP63JQ4aBmDqhIWGt4wviBdX3D9jLVz9+BLOTslw9HulSupnTz2IPyp272gv9Y
pUV/k5ug31gKX0qYuK8fwP/YUSfUIScidQw314+5nKWnU4HKDQye/rgf20rc52YI
GDP0qJTGWmxsA0j1hKAKlLTIxOR8yRWYQ2g1Ednj1haywANeBDJGs+XZOQJXXpMj
3f7dA9yGSLWngtFXjBUrJuzwMN6dvVN2CGUlGhuphGd2jL+RWGc8KasZ3+SdH5Fc
XqMv2FzZZnL21gzGDsC8l1nCmNC9e740U9ANhJC/wMdraERMm9W69eYowrNKe3Rf
nSD5U/Qlm53bP0JW002oAumDQiCzZGXhuT3LQ7ukYXhjzl6rfEWPRm70Xg0sw3x5
XTVlbP9yHy5ihQsStkC1j5zn7JUyJLlRDMI8yKKRNg1DvEuO9xbsHWwxSpri96VR
PQEhJeKyuPXbqv7QN4ftuTsi1FNAsAYZjDVcmBUmtX0K/vci349LlDEMRFs2iFl1
NjIfb0dOl/iIvp87ZM/ThAppTKJozltER8yihyKB0VIvXO3eIogZSrX70IwdEn0j
D4g5cYO5XfXQ64xYu65hkrVypNBpNTvCofa49RWVNhd1d9Qrx9cf95xKdqMblqWi
pMpjI6smFxF2RAz5POfG0Zo27twD1JjtfLJ4CK9aGdR9pTwohAyLHWQBmtC91Y4v
e81SQr9cRBiOUSSktWQ3F5iihjegYztH3Fuq0ooZfatI+/+VNCh6H6PDqt0lNpyA
9yetO5ongJwvG1PmnvukGKMEdgg8/Qz7YYAIiJ4oIl09vKeCTtuyJiesPn4cteZP
fuGHEygQlBjGbmAWgf/Kll7w3WAtpqjimWRc4ccD5bcrRb7q1DIfZkXl/+S59/Mh
O20yocO+cMUYMkpmf2fYiPFM2qW/1bV/OyXRGizUx6fk1hSYF1KCn94GNrLLT0oY
SwiVwWOEE5PmKPEUi3hUoJRlaY0yQSwMOHZtrXDs9ATLTQ2i4WEYpKOYmXxgUPF3
nSlzaU13zKRopeU57mjc1AKUNTNroeV/ketMR0OSsXYS1HRIDIbe9G0SFIYq90rT
MCO88N390l7lI4q4n+LKtRO6ZnC0kdyueozZhjOMXNqFo9gB5NpK5zebJ7KNvdii
7CJ8SsE6PaN9kvUtjUIe+dreuSEEQ0UQaT08keZqOfJ8/hK56jviO2hyFiVVNpbb
o+QW9IgIiZeAaKScdhbEV9Gp1+mJUZglBURJephTEChm9YJrmQY8kRGGSHD9fN+M
7/y51SNNPEDq8bKKRvka/ocz+0BadnT93Px0StFS2vGI+TxCkPC/XxTX7aNc1SbF
A72gUoOjgfHS/OKgfVN6jmDMNltkV0kFmny80WFSMi8lwI185uGdrp7Hk8CtoMso
qCupnRAELx/MvwKCwDJoOEpk2D/uj5pk+Mf4Q6wifnNh0Q2Nm2NREM5f96cMjGTS
aXTzYueti7L8+mkPIfs7VOFoDEJnLADKMqmYT3arO1BpVvXvD4Yo9o2kHjSUEvyy
Amfjo1PHeFDcm9BU+c6MprD43Z6DIywOmbam27b5sqCXIzJmruRb7booZEDljyTn
iqn/6R3CAM7IVxxs9Gj4o2f6MN3F6zRe/g8wtYYyaDqNZjnI6bz6ECN+flBEd0kM
tPPgEeqPgEArq86eqVAgbkhox7W90C1vmMHcgzql4nM6K237QvU5WgL6BRIdWgux
ZU0135DsKM0nNJQZgTR/EiIh3tsm5X7o3nGn0JVUFEQnpn1ARcFUJGcxTU/RwO7n
4F3jVYlaXV20R8XRdDT9d8HOOQdemVfwNQYfzdvGq7koGTr74eHWpoXblN5HXI41
I8vZmv5rfJehLa/zUV5KdM2w+SJuoQReNrckiRt6M81mpdjBQqyzjgWKiQZclnRD
thd/MdeLwAtq9AIW67Q/O2smyG2rxL1+aluCiDzcuLY4tTvMqQ2WLV9xsx759+6W
s1040OajGdMEE5Fk49GEjNDzJxvdY4H/wkSLPHW0/ETtIEg8XeRy1qrrkoWO/E/Y
1I2iZLa23cilUeTCLxtKut36aR4J0vbyMaa7DBwIcYaO6GmBfM3OP4sk/GYVFrLi
T/90Th5TekgVp5gD7i4/hVDJZ4K7V6Uq1q0A8EPm8u3qYW60Iop5gG/S1cwcwiQR
tN9f7GzxJpBgmpqRLIIyRhw5mrC+tFopgpXAoiMUFuXBhJ7oITHc4kWionVyLA4a
YA5tZWZEWzgL3UHTgTGfIfkk8di+8QopD0obOc8rqueoZMESegFSCzYv3N73mEok
lHoplSYzoIt9qjRN+cBrKG3mZYQxF+ubC2K9ZS559fTLKGiRXE7oAas9K4QjQDfd
v+Sjx1+VTU7oy0gdurOhMa0s7QGm0c7FDMaZXRW/BieEtN5AKYurix35XUnKlRCp
EZS19IjSpfTxe4d9V/Z8Jt+ZDIQAYGNvAfTzAQhZupqI8IG2ccrv9VlLdHa1S2NJ
Upnk8ZVpZi+dV9fKLsh3Dnp51FNWiB8Ba7HlCe3yyjMozXE55ulkDTngWv70z9lK
rFlOoiwZZfpft6Tk730G7l/ytn2ZZyGSfIlak+beK/jthxWUNtpuo79dQI9zbI9Q
w0PIct2uNxuFAfwfjAc0R0C/LtCB1apvR4u+dO1cOhBe8+Uzy67bm7W9+H4B8gIp
0bBgRhMZggDFkqw71SoOpz/1l2VwlKAPPqKA8gx5H9lOGrdmWj3I6oRb84apoOXK
gESMZy/ErGHMfWupNfFlep/413RTr0SYuMyAPM5xM+laPLlAHrAFJtEuTZwCqVbq
sahGRVktFtH+zi4D8Fqyvu+g2lUrB5HjKmii9iPnlangNIAazjWbZ/Opg34Ma257
jC+TOrnIHS/UXtjqtGDenkKuU69A/6kIPjEHpTRWtOsxyRkU5OeeLckVH+50TxAv
RmxQKiS8Qlceq9PEDifCi06LsOIXdolKwFFC9nQf+z45yTY1I0WQL3C49R++Q04v
qClAsxYfGFcKxYALT5YoCtZyXZbrh6xwmQ69vdADi3DxlUo6TMqiR3DVLERS7x+r
o3168FKLNje200pac8ESASdVZ9a1dvPnxd/D3cztcKX1qCyDD3JyFDx6RyjMleHk
VVoeJBKbkTLUtiyASF6LmR8HKfIBrj079X2QMPb6an2+uvDDZ7GZ/XVCBJ1Mu/vM
zonFAWw46dA+NF4Sv80yIQCBBzJKuYh7KM/kp680XVcL4bGdmj8yVD/mWaaN2yGF
vAR8uzDjoLJ+qQHG5bLxJvP2hrc8UK20MPQiXFoCFU6l62rY69qXlZtca8z46PXd
3xhrq8PRVaUcqvcrkY7kqx0uSvpGklZQFBV2nmwvxvOOFnDHYgeHsEclMMAjNc3g
pCWkeX0xsVbN27tKNNtdnDwQCpZ83mCwrY2MjJTyNxsmOkV1TtqeMxCFZGHIxvbm
/IeDOEXmfMb9VHzh3/G9fNgBRlZyao2OY9TQtQcxGTYr0O8w6P0Paj0PeWWyS5jj
7gvb+iDmVzT+mpHmm/R3wRXMG/F93eQ4atGVugTRV8cuxCSt/PV4uu0ouBo23oip
McrF9sVrcxOJ0lhbqBP7N/gtnrOF1phfI9Y41uNzuLI4gZJtVypTG0BbnwrvCXwK
rbsNcsnsYfzZzZNFA6UTO+ddeI+aN1nsv9UJJaW2c01EF7yRGIgwmo1iNClFR/P8
LD5Ps8DTEOsIHcHtpzJMvF/XbVKXk/h2P/dSI1WDPqacpwu6NcG8OjndNtVXHeyt
GI9kJd8SPFaBviPGiIerXTTU+gl+1ekLzDSr4mrA2WSZr6yweOQiCdqbmat2dce8
sF4cydewPZqb3kFN/YqjeP/pmOvUB21wI3QSBxq86mc+OtFbDuSxDtRRyC0slG0d
ngYOIx7nXBRqAcDbdoa32AmIV0mtSONgTSiC7TsRO5N7g9HQ7lO0UDRmTALBMkd7
ndVp3qbIXYgdrnJdVDffSyY4q0yr8xGuq/giafMLm8ttaQgQqN6G/bUdJ4An4rOi
zA1JQHfeUKYcybjlM3yxNIZsL7Unqvss2c4QD/OGJtzJIuB2OtiNk+Ue5PfVFcuK
MDg+D5KjJ8PITaXYrAohw3n+J35kfaTN65kIrNuq9TTfPmn+MOmEpfMtz9x3Fqn5
48xXpmqbD2oF53DEhdxL3OjcmX5Fwzj1VtWhi8uzwfsqO44fmV5UwQtbps2HjYIK
vgkj1qRDor6s5Dt2sZr46IJPGOvxlEAiwl+KDqhu0W39KBF2JOZ3xD8IdjHvRqPU
WoTCRbEZ6mUmtsnfhlNnwNDCzcfRyDBQM+E88ux2iN8ADwsusT5SGJKoUbV2p8F0
d9hF+7GHogcZpVv+lJy8kAYG8ubMljNQTg9WLWtDQsENcYUQ+TtdT3EhcfYZK20C
VWj6ADlbV1M610QECjGv5Q+tqWa/Vp7Y2uOIypGYKOUQJuymZpUw7gyfA8C/1i7J
E/XL4bJtglSI0xMpXPg8v+Frmm5AXYPlPZn1uyEXqh16xX0LKIt4lrxniJ1L8R4T
Y2yt0pV1QhhVXnG4DYAiOFgLAw2vc1gh7HSjUT6/XXrKliZG0HsD/r0fTb8hqhLk
W6HhUAQl+AzzL0VggSFKt17nDAkYNe0ip/fEbhEj0cLtG9xMwEmzZVGioqM/ft44
ddOFHImON0aTqBJ+qbkPbDmyx9z3mfKdk/bkgc6/KF96Hb2W3mFAAaY5NMaAeR0H
dn+QMyxwdha/MSSwCnNMjWwhCTSCnhrKl5p8t8Lh/KEZpjaXvYvmi7C3y3r7gTqB
1I5r3nM4hwCRNqblVx2sVhspWwR8u4o+3Je4LYcPum6rAfohgKZmkf79U1X7Sq0f
JZhfg7Y989bw3/uSBxaeRHLqNLa5TPQ+DbVIi8fi8w8KIIp8ypc6YAfDLHRw4Ha5
28a/coLzhrZu+hbVAfu3dBxuaREh8KUM43j/X79M+HMIJrT8m2u1H8EoFsJ7Q+Kr
AQhm6nCrsaDfw10RkxO3lCaAsVvzHm04TAAHvGI0/7HKAcdNg7MarMKw8Rv+X0bt
mHauUKfYmf+MZLODeZlozXb+CJ68GtnZtnmbCMaqnMu6cyUk23d+2MI7gd2c0Neo
Dg1TahV4SciwXMWga3/L45MmFsipx441qHSM+mv9DyOv2Ss8kIS3Kv4g8czwxp5T
9ZsczdnmOQs1794z+9jAZQLAC48mEr0ezOxr94SKbZlAECezxPAIp3y6PlF3TkS+
j2YX6lNYStpF+D8wKf/KXzEFVuOv9KKQ8IyIcLz6EV6TXtJwT/RUSfygwYpouQiZ
+GwWgksuJKSOxjamYtp3I1BZQv+v+CAJ31nVfy7qLVHNXWV1sUiXeoLHQpaKd8mi
+/dmCGzR4oN78crMaeih7oIRDxlhed8mnRbqQIABaCYm9oaggs5ixqwYQjaDwx9R
ZbLijNLCn+WRMUi4RdjAEp6sO+K/8T1FvlmpyCM2GBBLYHdbKOO5tAc3Rj8JwdFw
uQo1N0dXwreYR56ahNYr4tqwB7NKeJc+j9PuPpauwfj3jHZW1GziXmcyD4vsuzJ7
idW3NVgMhCu+eEU8RRqmXJ/7QbZ+0+HYrglp2M8bGtfPAUuITFoMwMsgcIg1au1W
ufc7bHEybgXZ4GCM04S5zgKft6FO3Guk+C/yEeC2cGNwL9yQB3QKH1fDk1Xd9ksT
OxDOxNJyqgom52ETvh5YiYFIPDcT22WxYOfYL0aI1CtWPU7YKWgCwVjpxGSuFZaK
RYP8Z7Bv5paxYJLj4cfysSf8MSMMGv1a7UETCVno7TQbOfUPBekJWonGKWErtg6n
JueE3Bn9EuQNfSwtLrz7aDWeD1euWXPrfoU2ABDRJOojccnt9zhK20+nCPsa6LVw
7hLranZ2CpxF2WxnBscSfTcrypyvfCll82Pigl7mbQCmhAy0FHgAR+2dXeU9Uv11
Jdcj1UT65w33n1TIYYiNGJfGZXr8ih3eWQ3Fj26sFj5l4QabMACV0NuKR4FUaxKr
3QwFqCm1G2N2Acwql5kTwdmP2ES03y0cZ51FttfMq1WqXOT7qgva9q6ZxUkGCdSY
Z01zIyUaRuDhCSDcJjVhCgRUiQu+ModE6keO+dwERyWH2GJbbkOwF4FwOcbABkiJ
LCagrdgyD0zuORuGOyBfyCeolBcV0+6mRmxUbeLtGwXMMjvxg4Ybh7o8lOnMBqoP
QeNfRE7w5Efi3myLqpjUirRpScG7Y231pKZpGeK7yN32eC43yXAgE6fBCJjYzwO6
2kiLYU00Hm3YsOlsPUqcG6ZMaEJWa7uZJ+IUarGjszXHZbGLB+r2a3AUVIzID9g2
RgLZkvURMAJ9CwCkb+UKFO2okGavxoLbybHu4uWDQz0fJd2IDbJdMXJJJ5I90Io+
VSOvPlT/Av/771MpoJ7efAss9KLmVemYj0iszRyw5wasV4oEHnMim8878beONfIc
5OFbM7ZABsDl8gF91aHqlVStGQASq3S3b6nEx1ycsOpoISnLpJA3OUryXPCbRqcF
1Ll0lQmFjT+wWXLJpGrD4StO5F0cbMp2mIuGDS/xN8aoIxSQLCmUrQ73Iz5kM9FA
nhUJpjVl1X/GxM++80y9tW8mWFJSswidWRTwM/d7royZWefTlcloINrff5Kn1Tct
dV2rq9LzIcGUoo6wDqY6voVBIV8PfXW16GGGQSn0rzeW6g+ZoeCT4DJRHrl1qHaz
kWQA9x3GkViUPL6fvfkKBV8tGUccHZ64RHqi2xnM4DWw5IAEFngz+Du2nuMxJKfV
rm0bZYMaszLs9ORtsiAVkHPyt8Js/kVfU3TifovTXSwCOi516nNaTw1N8sx0SBL4
6Rew6q1d9tw5qVER7wwZszxEfsV5Qmr+kdh/bUGjkQahQQW/PKPN4eMqlUgj6IXp
jbMldIf9Zz13alGGLkA3xGd/qbshjp2boyyvJ5qjOOhH68UZr3vUJJBCUFounMii
dDczwyJHr4qMVW+2TshRGv9Mb1B7MC8zz8uzEMIOY3XsyY+VCTLftVTzec/gxi8g
kKPvK43njvj3AxkxznsF/tdn1AGMIDlAsUYKHQw/sX6UX12lsGH3LYZhxuiWqnFV
z6PK8Pk4MR8o76Khqrv8UGSOEo2EggSMbuQ5+ikhwYlOgStmYTJlD5+NAWzuB74S
Dfh2EPH6vb2ew86AczUTkZ48FlGpX4JZhRmfklGAl44kbPeAR6YSuckh00R5gUWL
jE5Wd5QHKJ80JQ1ZmM2tvM2nPNFHXa4pZ2GlEjo7i1Z3NJRnkacGLK5hzZEe7QpV
mUUIiZEVxUoiJkFiu1KNKYBOURnUigiIDhOdPqLha6k/nK3rkMeIOh0xu487cmFQ
M2n7MAK3bUHuNqcAKuyDzON+zWkvyXjNGTs+UJWhrmkKvgmVUTi4qZtZNlNJPpEA
eHIeBhkrbZOIafrijuwYQ8zuoCWRmMXxXS/DGBAr/pvh5UItOmFO69RFcUMO3ju4
b5N028UqlAc0mJkq9sMkAotnenpFADj/b+03Z3TQpA8YtIPfj33I028FHCj89tVu
yzPURVxbT6+lcRE4DQh8HFeyK8oyVNOjsGH8s++DOM1/yfqYQIFqT40+hYSJch/g
zPvO/JONVfNkkRrMaaSPSvfS6NFQ7ysanfjiWE5yL9FFzY8mqluvIyQpQjOe/Zo6
Kll0OJM8pJF8WZVydYoctYAmv1MWn6UG6HC/aiyxxlJIKrVHp1T3pVWYrAWCDN1w
hwVW3zyjv85Zs5N9xqQexqzEkD+H35BLEHsKOstP+Htu2L+fdhVWhN8tkcYs2qpQ
yVMHKPLeIah5NxrUyUI3JXKdKBYISUdN0pCN7wqhN0vuAp6HtrQ+PmBVtUj55h9W
Zmlpg9JlxR+tldVAFj1LCEKotm2eqFSMXyebdgh3y5LaLn1tHDE50o+TJFfW2mP4
nrSNsi7ag2CvSSDv5IDpa/cMLJ9Y5BMrYWcUxHfV96QsFVNqaRoHu1ZD2jogKNvT
mmaVQ0i8kSkDE17m+UnffFB4peI5LvmHBqWoAjHnG/03w/G/YR8BihbM35HDnB13
wNLlDv14oJcTUE1CAjBU7EH3vOdVLQS/ayT07nWLEYCoXaWx9CqA5ihj/ZIIb4FK
tG9du3Ao0qMYwS9MEZ9ObxD4VnoJVTeWLeHRRcFsPk9ixiPZcpbXopG6ImjPfEAr
Vz0QPqSQDGNzSgZg0ggySKHTNrxDS2XmGEq+Ezc964T061ZL5PR5Jla+tirKza10
1B/qILXD7xPXtWhQgej/KmyUGTwteHrCoAsfp5rrcdxSae4jaxYOdZWMmUe4xR9U
qE+EaoGZZ9rMlKhRt/z4g2AKX36N1OHSVH3QcPOlZNDVifSFCgEjoh/7h3UNt7rX
0wm1V+SI2WMW7qLfuYmu8oQVHxQ16pYPFjtrdjioV2A+Hvd2b9SpLA8tAZ95g6fp
+x4aj1yRAyW6iIFcQbL/aPoXT4aMaluGRGlor7CyNtASud+2leZTcFJTccvTPM9n
oqa0Df7qx/ON5oJTDo5H1i4AOTboq+qJBKKY5RON7WfjmZ507Fyj3WEttZsGLqll
eJBA1p3YojSd9lWFA+xDIpRCn2wAb3XW9dnflw/3onEri4+AEkuuxGDg+Q2S3vFx
jwPgFjmckjxWV0nIDvmQ/x/T6SoiKyQLPIH2u2hIRPdBIuWCdvQJoicIXg6EVsUr
nEG9u1mGRdKRXN9Ag5jTFwV+PjqHuczUCD6hkzBWrX1RxE0O3Kiysn6zd0gDM9Ky
FeCVZAZ0fa5aUZotVRaY2Ln0hUeL0bauGa846y+qobP1QvpMX1z7EXvyQwRhYg9t
75o+Y106uDBVOjmaHBeGwQJ5VXxLOHtMxvuW5zB3JVRTxgH2y3R7dlci4ymcFUvI
pbPrsqdh8EmQb8HeRc45rA1TdYZDKsi7Z+u7DZ88Nx4ADpi7qrvCbtxVy9it/lr+
MbKhUsPQnVBqjLSVYd2iwZYlEXXflbZEyP8I9PgjnCIPb/80PBag5YYQxbIqVK6q
jOmkgsH8wmyVaLkwIGUE2fhuTAXrIIJZjNE7P3IPHZJ26Jr1IbM2In5oBMgFmXrj
XC8iYxJuggwpbO6u1k+kIPpCIQVL1QDswyEnGogNVsimkPbXVwqO8lL0i4sBhNgv
hkywUdbVTb2M7I24CvqFjTQXs+rrITqB5HnhiD2ekqDVKUDTJPEhg5iTtQeTufiP
PXY7EsssFGtggRZzP1VuL2/2yp1UR30WSjFxl9rEG4dYAySouI5szKYPAZg0xMKX
lIKvRxWbx6d+yUY8uuf+ABrmmT2wlJi2ROqE8wbwOrN+CHSB3ywqUuTAZcRL6NS0
9x3cpw7ZTaMSr7qluIY+y0Olj52cLysVkeqBmmJ7s109Q+gOpPh+VPJ//MxjC8j2
dXZFyFRxZ4F6u1U4iU4zkEMZIEn97QLMSi/m97/Zrhnqag6e1T6NzmDhn7acjIt0
CV3bX4fHm3lYqncAzFVDQW+wQXR7jRU8994kAK2AIfcto1uGDqRaa3PpKZR4TO2m
A2eFE+B7yjueMs+51lfjWJmyQr/T6kfy2de1bFuEhUeG6EQsrsDCle5u1c0h9Vm/
RuITFWYouOp/KQeqzOBWZGut3g0+ddvTsCByZrTa7nuKW4BfJz+hFFIzKVWrEuTa
9x3wt/N8Z4uMTNThkphHNxiKvDLe4eSF+Q1xxZX+cIIjga3szBF33VpkI8ALCCkt
t+vGmjUhe7UPBxiUV8/ioWP6xZO8cX2JYM9OnGSVMPEa9fe5o2uiz6bGgd7/VwgI
FXc+nA+NAcH3YR4M8oAg+ZFk4f+B6LpSZibNeBMTVIjVNr3TW3Bj6VqsSVClxIOe
qoppY6MUfjWJQd3x2TLX0kGs+i/2avI21/U+y1uTWv34HHWZnA7BpGtp+7/wnJnp
J6r/frJ+GyC4LepS2yHYdLx7Z8IPk4cTBZKQEw/1aJ5KsX1wiJUWU7mnltMUyFTA
PXgBdSAHC3aJYzm0NnHCN+QBOMjpcPTYPfmJBBkijd01/17HaERPppCDBZQq+YWz
nfFsMX7Q72WpfvJEsRmu5R6pHgB3lFlKxFX/53GnUPNld1rvnKj6QP3HW8RJWfUI
oIdDyCHIMorvwCVOvGaQQ3Rd+kCOPirCLu60Jx7jRVV5+/YWN5EcPveSbGcbifL9
xGg5HVy+Yp4a7XsW6jJAHhxITttKnI4O7z+cjEdq8vq3q+jz/SaEYSpXRSDBTLSv
rjqRLBwSUIK1NO9o+USd9EYFF1JWcZmBnIBEtorN1jn03wlAEj32I048ScffgD+z
rIGIRTY6bDCYYea787hxPsrvCyAMwXY2AkT646+lRn64yRqfYln2/O6wQ4wgk02U
C8R3RS3jbbT3kO/2OkPqfl3XOzPN6fpHS96nDasYRKpgoouauARloOkRil3FCnto
oKAxxMgAyMRqwiRdWSjGX5Mhl4Facd8sIl1FA2feQbZV8iSNclPKGDu3oihX5luU
2UAqb3k+2o29Pd0eBbxmBT7MUe0XTRu9eS15Qms+BK0Oemj/7eKY/BE5vdqZPWDt
MThd/iurTo+qRi2iAbguk/o8jP0tKiRLXvlLcecXdjBKh3DmpVISPU2pJ5RYX13B
uksZnrpkq4fRdK25pluvoH5ptgLNT/gulIIU+SFFr7QP7MHS+L1KYQFIoSXeGapj
mraRqrdz0G6HWpiT6iy5aYdRIcRSShy83tQtNqvdlQcOQLkeLnM7m1a+i825DD0c
XrqXesW/YlL5OxUrrhUFIGy0kGe1LswojGrGdI1LBBpLMQv3SQ6H9mpEufqaLLfN
PrP+RN+DOmD67aJcB26w614N+icLqgOvALcSqF10GTh57kuPZ5hPHNFeipWmD1zv
HOnSO5/rwA1dk7ZPHMTpSpx5US/I73tOGfqegn2ObSfhiJEanfSIDrZgTVjXnrih
pZp19HbJpYfFEs8TyTc3bbrVqFyGGBbkK6k7jDbH2rjt1zjBWTriY3VF88as2exT
c67A1c4IUwl3TVT/tV8JmXxNztrHZeIEo+J1iDFiD8tD9Gp6K1vslzs+47UB0TK5
SXhn1iHtaEL0oDfmCIqRXn+Vt1uNknJhGYRVoQHVVWPtOmR+eF59Czn01J168wZo
eNWwT+FXtULh+/VEwsjRcaPY21SgHKfSKyR+DMPxJo7l8fuiEOCeQeOY3MPiUOBR
Ivm0MXEjMtnOrDnDGtMCNnhy3XYzZeOy5qgjPEruvH3unDd0ddSR+wfDmM7AJ6Hm
FTg85gpWSBnpyPwtJ7H9MPW3+mgsue7+8RKyEepXeRafKy5TZlXwlaw/xG0utHnN
Nd9Xqeg0rKbKSADbRm6nVpYH3KgQ32OQEnrRZfEgAeM+bAMhztPOhXSwGw2TVPer
Z+y7RGrzuXBMwlCYxv5Dxq330XoqSoAx+6PkVyoLke/Stg8LAzp+cVWqOJ7T2GUC
DEoRUC303Si36kmG6hOVxx9zes05SmqkxhJQbn9zx3Ve0A+U8w33aDptoPD/xdx+
YCHJ1pw58fteUMcNUMi1hvykZb6WbmltC3bwjihj+nZ62r++x7ygfxAH0TM07w/4
AnD9E8kAONN+5C32cMoVEb9G6oJK62czfC58rqxlTsVghV3IYsV1m6uoApYHtTRG
/i7ZC753LSxKbW6DOS7lu5EmfdSSf5mVeyRc/r6Ka6oOn3KHQq0fk8O/3NilCpI6
RetSRMp/pMTlXVIgDhlZwOgPVeAs4hIR7p5O4TxaPdZ9Y61ngVl6DrFZlZ6YHkUI
P3FMtsHVeSaTbIPSZt1H0K9Cbu+X74tCGbpgcVDuDaILZp2/EqzCkEUydlizmIB3
p0MgEBq25Mm7cmWQxC7FS3Y4Sfazg73isrR7iAmYmyTVttO0Ww3hHT3QmHZhQODp
1juKHNEFYswtluH02W9Agttk1+6XVugCg2ElS5063CSfFlNXg4ryiAM3GtxdykeI
DGADlnctvZWs5uPzUF/PSi6U6SwfS6xKS/NZIb7cXNpap+TU80+xOeNaxxzSEiBm
Q3uFrcx0pWoPvhHgpz+XrdZiMTjqwGULr+H8vtcKElodUczaU7lUOl53CdiStREp
B2/jUtyE+5lWRjbh73BId5WgulBUq9cPjZuPqPJdpSTaM77Y9scpB99kM8gAGmzM
9nKmBk8h4KcmCfPrTjld7UamtzO+Cz7if8hIxSTsMTTY5+EwtxQiDRAQ1Isiw+MT
tPKiYBIM+OwSL6e0pzHxQQm9r+vVMa5dbS8i241zkfqxnJTi5cmqTZCPNiKfd2iz
+j/iHGZFDnw9mVcmbB0MUxVOlaZDklO8eZ+T6uK5yNMeUVbcKJs/eK4WbBZ0+zbl
tfS8c3kZlRdTF3Zd+iJlD42AVljzboWfe3r7f3ryRVmH4ADe5k44se37/sLIlUik
OVPikKs8tdc+gAESKaqtHAsAnYkG8CFaO6l9VW6wsxuiYbqZ4H62w0vsgHLVnwSn
gGYHIJZiPgQcYg2BcLxtu0fJVv+peeAJh1d6jXmpm4MKWG2sqNXYQ/bL+3WBkqNr
H9fsqMeg7vUBixIW+EAjIiNkBVIDMtdJAnNsWhVm08iezPRyk+yMoa3pmE3Z9OgT
GuAptFK9IE2/gIwz/vBDj4tagZI9O+qIPWIn0LfO/hQRZJ4IzhFnNE/HyzlPzGz0
EgVBnaX7P9kYMMQv8H+7hRNKoVH3K7MitP5hU3h9WuI+gp6XRM/OCnxiE8aKsoux
WllK8O2Shnu15MJ3RVnSzS4kNanTGWjQgpk+8M8fbREiOhisfpcbdVJg/ppmpqwk
FF197T2hYl2LMGrpi2PmjPdqS3vBeAvoUTeRwJk/iZGAU21BVbuoonhwOkstM9HM
nCiYytvKlqHzXO7Dz66Yzm1hZY4KrY7m3a5qq++p/lC46paKjxIaIoOthxZYHAx3
s/QKOcfF5wAdy66cwqWCaX+QSExziRfyTmPdIOXf2AQyUt4HKaGzzKXW5yQP0Nqi
x2rbTNMKbWBceggTE0aCziksNd7DFN7yX+ORafXSMoSPDD6myJjtL4N0JGVpBfK8
GfxtT2LFPDN9VMnmTilnBhaJBn6/6yMzXfRSTD3yX6Ne+9ASy3OWY5r+FbqfepHQ
JxYeEBDIvm1HQYXEF3QIS2sUAjTPrvBx73I7aLiWobIVMsVW+iAHIOqOQGUu0dA4
LjHKB5BZfBmi85ccW1EOgRvhBiWs9FmWr34UIafwFs/McVIFQuTBWCye+/f7Ddoh
XP7gXIsIbZX4Yqs6ac6Js/E6IKmC6hxd2m44xOnBue5XicJSG7gXsz2qIsCTKPT2
eetk92tX3mTfo/ZiPZB+YDOmfRAaFhkLtjdpn7GQK4xy6c6GWerS73umEHHOUX1h
/wL0xrumC4f1IUrmhIO86KrkMXY7d1BVW/bMLX8mDksg7PTWOxZu7Honiz8NYDhm
95HmikG3rTiXuIOCAYEA/Rz/L0kZQWNZEl/AQ8UFj37WoWMnfyNQLc746fr/36BN
xVSASMYaT2X9uqJtcjThcUSj7JKn4aSuMxdduCaNfzdJOyVh6lRBV4THc3HkgXog
yqe63l0ugD8WHq6mfmz7mYC/xs3N/X4Xx+f1kR24btI9PibucQAEUiMDW5qq/fs7
cNeqm7+Mcq5v2rXSee6WfhCGvU1KXwDsTvFnLfkYe9umWsLJiJLX39A1GYDL+UV/
JocQT80BG5JBvJ1UC05ZsLEOEE8o6NybYbxLjGTEo6SlYN+dh4YWxa5buXLYCNRJ
+TVZmH4LLRbkQdPH2iYxElQVo01icZsSKoIxxe0+GfvYwCjazrAG+3oLeYn7uxPq
Cd8UajmQojrMPw8OSNND5qbNHuanAuQhLA5rL1OvRSkgPmkI6p90NWRx1iREb9fb
k3EWZa3VMMy0fO/FPc3pceTRNXMDLaJBFkXDMLGFjcj3BubSpodxlseAzhlZdwN/
PEwLEypQeHEMJ7ou9UbrtxKAAQNQGHJYXBWcwqEDBYEPtyTfojEGqGRPqBMIPQnb
fTjKO934M9csmUDFS2lBRrPY6/FAvGI+X4W3lyE69PplNqtcyMhak+xadK1jICtj
ODYM4bL5ZnsdIPyjUImLrdRUonNC5UfdOM/lPwqb5Riiq8P8VKw3wgNQZLR0YCmd
YLND7//fS9SqsBmCIVNn73xe4EqL8sH3iyjPHvbZrdfZAwjGp31DZ4L+5YvUVZzY
GdeLp21YAOZEAMGJVVfcvrCAvOMcfPHW7PFC1rJ5dVuLu7EcCjhTp7zMGtfno6na
vCHArVRF2514oXSSYdl1cNin0Mij9DsrjkKyqWkpqbrlRNZYTfBWyG4+tFx7CTQv
yuUkvPyEEMVLMnXNGszXg1MhR5zozo7lqX5f1toB+tWP8Yl/zzN2hsbURHUM/KaV
fWxFHEX+Xr1ZdKg9JKfptDtUbfyse3lBNb770/lXMwyYTsGWocjWcsXa7z2YlxFV
WAFUp0AYjypFsDdIodXhcpLaKdUTyjFT9dQrtp3suXECHlUAw6HzNXvJbbPSbHzI
zQ2UjMyX6hV7M/cV4cQR7pmpIcwwjyJijkObnszrNyH9121Ce+XFec5ukebscRGr
uEqFwlryWgnfOm2PPwC37ofNN7ldEnnLu1DYj+aPFo2mzDw8UjfOLIVyH82WwmMG
Ws8h9kidnRIpgydyTa5UDBaEFnzqWNmuYD4jmNO38YXtPAMWprSSMeOM5q7YI1C5
8d/Gd5h82oYg89ULhD81sG+Boy1Bgp2vp2dDn8O3gZR0VKKlRf5VPuqKMhV5wUlz
OPkhIi91F5hZ1bO0oMmbdEEJoQA7yLwQWDAMD9PyCEsrAtEsuqRbXdMBOzQVOQ9h
qNxdHnPuE7LV5oJwUg8Dsm1oCjwEzSeV7fh79aSwiksc17xNjEtCSNB8cCaJSpBq
1hJlZvc5sQfvrKJyL0czxUWtozig8A+kx1HMh9KBUHWZ59Rt1T3LwBW0mdQzNBIz
pBySBtxCLy7NmpLxDKwuePcwQAMmZkOZnqRaWepqiujncQ9kjzC+QL1UU9/yxDIn
X6Ru8Q+PoLXAy/d8NpSFh6JT2AxqjeXBLibiMLz1pkkGwQj3Px7pxLp8TfJ83zo5
9haICscBB0qB/lcrP6tBIxAqP5wAY7QJUck8O6EkFpqKFK0/Y6zM9FSATcdgiZlJ
k9MN9L+62XcrWEg5kmmkZZC+fzP+M5dC3g8J8DQVoe5r1N6teWG+0XSgJkyZ6cKT
doabv+zipNE20bl4/X0/YII440fm0YLFzL9iP4dWAHXK7Oa6ymuS2I0C3ZJazKSJ
T6rWhlSdI/U3i45zvGzkBajHjlzzHQuCWP4eCjf4GCXt4klqH3oTrpjnMmfndttu
zHGHlNOi0InGs/B0DDf9dq7oeYjvHXt0O1IsX6+k32Gd0oc/U28+prqShtdiZuAX
z6K75BV+IsmkPc0BPXuEGpZS9BZk52Aks8EIjfyM1AcDS9LMTT3clEvWgDv+MsC9
mHfd89xzSrgTSBNd623ub3d9toriuxD6apr7QHO5B3BzOydOUDkcYxecGB1QLbjL
3NAceTqAwW787ilYleA9WWBXuVmBMY7/tvjr1ubmAVzJSPDSfXI2SuUwqHt9Sca2
EpoSYQ+yiny6ZVEac9usF85aX/kMi3Ztz4jlUUkL7GIpyvq+Tna1bMsbHbqRoFNy
s45reSNScaQImoG/Bp4FAhR89yRo0hQUGaZAoYi4sfsvnOato1d6akPDrRrdidKB
pi/V8he8tp88jaL1kUruUADdjfNETXiDy3i7Ac0PbedqVbumCDOCTMc3by/WTssu
R7UFZzHca/9g6g9iYFflXvpbjfREuObXc8wYEzw82Wc/FCLbw230Byr4KLsbjdjP
Kczn4I3I2pQ7InZhlfUE98MA+jx4eDmluE7M+dBtj+RcCBQw0OOgJwTqQGOjM0Th
atq5Jjg86FNreLoNkz9NiXHIACGK3fcci7QAJBbPgV0OQbx+AcuR4DxsR61CZldJ
pFiNxy5c5ISwNgkreLVcwjrTLkM82D4C/YjjkrUyjdlMeCKxJgU0shTkzpOGeaoy
SxAXe+oZ1w+SaUEL1P9/Nrfi8XCJWkvA6AzwVZWk8JcLh+5Zsm/KskWBM32jjruQ
eMg1517wWIqc57NFPnJRtA1SqHiyJi9vj/aIavuXGYUzXQyhOFfjUr/Dl8rRVjQq
htF03lwYPGyyvdINz4+wOUXy7F1Bb0ai8zbS2QHmUEIKxJT9lCv9DQTd8tTYoTwb
5RaF0dg+La7WbuUZljndlqg8SUsDkk63xwTy4ASLjYyNiEzO+tRtPYp34I9houlB
CUsLku56egx8OENGnUud3c0l2u3nDHNvJTMEkbgjiEKA3natSZE1xvbfDMZ4OClu
uEyDYjxPPZpCleZchl5voGSoX/S33aN7kVh0qCVr54m5g24GeWNhKCOZtmlGLllS
ty7DOot27EWBisDYDeaXp0LSkgLC6JV+gOwtCEj1XKs93SNO+qdfH36ody6M+01S
tvL704HyABSQPfOHvONsgIkfCozH/Lq0VZM2YVDQ5lTPEgM64Xgf1g//SDgjSiLL
H+RetsmXSBZGMBnrMh77G/YEsMSQBKIlLzd2p3MSMlRjyEnljcAXWaLX25blt31B
0tYTf4yr9doI34IdM2I7xmglmtlVJFJmrUco065mXdk9Yx5lDSggAz+Vgv4lvUvV
dYat41Sa02lxUeFmDMEP4hH0cReB7y7YaForMQ5AyE7nfeuuNYaiN2w+gBTzojhp
8EJcL1AlKMZOoC82fRkNzkKsMoqzInL3OeGkqo4hUYMV24nLiCu+JJlaewCbBDJp
sSI1ILIcabpSw4j9jo0WIcTZG/B17+uNecR5zFJMr7QxBLqj9y8/eWvXv8aRA2y4
R3zgEaxDwBEKeWfCBmhqCOaLaSfDMq2dufT4SMbM1/tV0y3SyOsDd6Oy2t9UGtMS
rU+10z6rXhAvpXsLyySuhe5pPEcgz2Lcd7xFBq/h5FqOYqGoLIKTpZHJJ0EDQ95i
Cvwh8lSN4Dr8PhqC7i2xrOS9zGYZHYPftsHIlbJzT3cL1KSO9RlXWkohc6b+ZEEj
uzkxE7DJP0fDYdSnGoPVbPp9x6bfxH7BLLXKomJg63z+SPJ9l0NqRyVfXlolh37V
PiuqBFSmndjjug7k8FbefL26q9ddVhs/b/5oLWBY2qNg6AYLJhQDH1bPyXmeRBWJ
KSthMaOoWicilD4fXuQfIZwjXlJj6AzTnmE7LI+hqWD8gWkU2JCleA6U6kh6O7kd
9XUovISzzhkY1964J2mHB2QKO9gyv3mRFiNunSTDPHX02qmai+MZUnjC6ygyEoRX
aTn7dfQ6xUtEgAZ2T47cKFiYapxLlJBj9w3ugNqa+zLk7uogbviDYzMzTLf15wxL
3C1e+k1yrE+/3I3rPK3yXrnxHdAuZ/wMl3n1mmO4iTFsiR66Y+2BFm85DEBPo9Po
GuNWapqo8MYxpr6jIsGXqjZy9x5OhvhH0XFhTC/ip5UradrYl0dQIcJerfgxDfkE
JY7wcKNsofjzTwsUKnghktGlBFdzwz9vPxSxb3NlI6x6dIHLBlTXiVZ6Wr2Mw2Uy
bb6aHnasS6vkZXRMtWrVPKGPsonZ5AjQcQLoPUPEF8FuAa64INiAxhzSkmoODU6G
0nX73ABltdPirTCqQFvnwRKfuvoXADN2TRFccfo0WCFt2EYmYRd6+0RshYbWGEAc
O1hljn+VUCUF2xo2ishrZoFfyiMby32gq+jHAWJl3GCqOz3mb6yWMvYLGGXrakKc
TOPG/VSKNGQJnlQ376LOVrOY9kLtbFbdn1T464vT0Uf6M1YiEODAKxxwBNsWhykU
t72sj7/1r10F+fX0D7yfQ1lPE5fF9p9sgTrB0f+Y9AaYVKF/lX2+edAXYGg9fNXN
oCdbjjbhRSD1jpvvXpceYEqeqZcKheA8rOOdUKk8hbQuufFjOPs8LUMYJ4D4dgOa
zyswvqQmt9KcQdQYJQ79US4/LHz2uTL7A85y/kHYTtatPKuYyuGOEEZKmSKJ2rQe
pF/ehlC+16pheP3YsqtkxbWVzFHXF5qyJvW19tECJEKqTrbllr0YV6/+7fir77zM
1Gkfv1B+7iDAoxpW8OD+0c5r9sOLc6uW9KM22kf0RdSNDDLsn7NjOSy5+mgW2l6F
kGjJRyriDCvkMaIrf+0cEGrytxwulILPJ9sHJ8pSbNmRqZ4ZrX1l95PCiJvS49bC
TMY+Uh9Ll2ap9vyZ9bzb3QClG/A1PsyoL/y8kDkKF3lPR7sGrWIwilT+VXJXM3pc
i60gZ9d4wuPAui2dlvp8Lrw/iR8MKSR8nIWo2MfVfrL5jhaU234CuKZHVzpWMNdG
d54sumV+VY5n4Ff96vITWUlIS8K0zGw6+78PtgWP9hSHCDHQH6CbE1Y2iiixqLwK
hK62oMk/KgORUwb60PFScrgjx6tmdP6FMeplhzV2dbg909rZRJ8TWQlFkmrFjbUS
2ID8CfadNUOU//Cua/slLvGEpH48lmrvzjyj/RPTjR8gTFtN7bMEBk0NPWUT1wKd
jv+8uzg/2ybrcBfofKe5spMCHbPKaCLl+eKGsjH/L0KrS5tNaX7EaKQ1Pxm0mewP
8kvrXY79TEXEjGrm+Tz0kBeR2LVUo7p4txnik0nutvSbdrz/fB3Cl9FSeKqajKQT
Dth4Kt6Ui+g8L/Gb6qIGqatBSjwzAPZP1ImchJMXW7JE1LC/oMjvJzkYCeDFP1EG
b8nOWauP6v7u5Em7aX2c6W1qfNVnRWwR+EWrn8ELx4JnXAQJAiwasoq27Iv2VLob
o9McwoUnO3c/P6u9FSWDlbacJtvOMHuU1ZHSvrXKJOjVb1G7w9Le1mwS5wNiboFK
zGHE1der+4pQAmiX+05CDPFqigB79AHobwvEimNNk9LaNfVdLQWIz+EaJJrvJcky
9GNBf9+eSNjYLQjsAbVkeJ+AcFbJ5s5tPDeGW5nJSY6nyIzIdvztTJjuTFBXq7oy
qjf3vzNeOgu1OORWxq0PLAkO2KksMuGKXlVIXR3YtxBBDvrY2UN53pBHdTvrhGmn
kbPcLOwNulaLgQoJP33qg5n4d/InhjTLBcm7njlxrBvnlSsefaN8t+bbeaHUmtfK
wqwY/s4VEoGNtThX6bkeVJY3I7j/WHA8IGw5StZJ5NzlhjzfWiBRyqPWpX6tgl8V
SbwhJeImVF6jUrDdZtzirpXpXbz27euSdzkeY6cavGPNeIH7KgV9ETmDFp3bxJH4
s22g17kxWxJeQCzcYXvFzZTzEslwKBYcNWJsNwP0YM5dpsy5qrLP2uKMf5Qn2jB0
45KGLBuaFtz54lEP4bvtmkv3BkmYzMRQkcSUlgUKcNcYGPHqHyzZW7ELhX3xwdcn
ibH8+i3DcDuYxUEWAR0fk1IyEqdjTD/kFtYpu5UCq6N5PTE7M81MeHNCRxJs69ie
7isyNCvFLpAZsruXO4Y5YcKtPp17oHJaObduybSeDIvAjCY9Y+8qHfbRkkRfNqvu
1eM64PhMe/kXhMlTle0r6RQ6RTWew3Kw9sZ2dX8NL+M2VuivpWdrLok6EFi+VVUv
haKgcZ6t+PRk2lrfhuUGxZgRGtoV57y6Dc0a9C1DcKMGRVVO3WAIq+MzXxi648RX
DHzD/sV+z8LYteVo3Kx5TwpVRr1sW4oPQHOro3s6MzVC+u2OV4FMejkOrwCCt/A4
FqyQ0pA48rHsG9Ko0TBj+T7b+YFu1rBz9ssh0sTYDf3zRzm+HZZtXlmuu4wdGz0r
XXdVpY2qe90FxjG3ywYdxaTI7cosj60CibnB+PPZ1pbIpKA8UMpzAkZslbFRq2gd
uQ4s4XcEUPFI+tWxMW2B9KZ1t+igXeyOE7/qaK1rxr2SWS2LPPeMflngr/QMXxG4
cCdGRe2sWYn+uhATgSx53avqnyMWaY/B9y9EXHAqhRjJcS8f0BIEuBAXQ4bbVEyU
TH+D6pfqvBKdeVMYIVmoAHU0xycwgdAdwYUwbD2oAiS0TuJiYmUnaC2zt57332gx
6VYZa8GoD0dkG2qNdBvhuHV8dsDfYGck2yNKhboBPQCFZE98A6F40ggwp/BdDCHy
6Zulldvi19j085K35jMJAaj0AFexklJ13mko8P+w29RjwYvZo9PqR3D0e1EZDxfF
YL67L6e3z2KN33RQUEL1UjW7mCe10AeBaaGHbdteQIdWCP+GV5J96Pi4wIqfh9/I
AMQWgY76wch18d5EvSuITpQwABMd+2VNQPoZzQ7wWAMuo1phYQlVMIud8Sc2+lhd
Yho3zofuWuErsxt/zXTlOhJB8ZAb2Lynx1ow5g7hB4hmGrkPKAiHeBQPKgoCZg6F
hSsXZ96JQ9LaajL4yXvjP7rxdZ7p0U2zJDO03TOv6HDflh2f9f988ym7PAe7/9Ac
bM21S/6KAT7XdPTm2sim2sd9VAFGxaQ8lELFglRRdRnMEGv8UjPsh++7KHqbjbu0
w6cEBaDC5xwakdxzkDKxuAgUSzbSIy9L/FCLOW8aA9jDsmvPxseQWvI+NeyWnKSE
Saufhi54aiA3/VWOIin9qHUY51loy7La3a1E5oWFSg4wcEoc25v4hPX22c+9VTeH
NuirmeaVC4uFIdBn9xLj8Cm62Ie2ScdrTMag0OA8ACsjGWb0feP11ulqWg7W87kG
dxzQS8sWaMjNDcj/EXrKi7pCOQ97VOZ6sPtOYbRme0oFDvL0KIocvjfUBITNix+r
H+BTsZSTTAZ9KFbJIjfc5WD4/n68fBV0czNWC+1h6q5Uqc+SAtwuxQk6FCpkKXMR
BHeXezwVXFdLt5UeNwNTsD2qsOsYWVfrLKa4gZQIktcfbn/VCfHftlCsiw3KxLmJ
1bBqmnBir37i+vX6YsIR8VE+TzBcZc0VQMAwxGvwFIuL/AGycAKHLZVrGXgWTNp/
SrHb+tBQW6rk370Ld4iAT+DKrrcnBkn5ppJAqOO5OGeu5ThPaXaJ5v1ZUYO5D3Kc
XS+wPHAZb/eZI28FbMh0VmBLnBiGwUKV0N64AaCcVKFJWM4lQ2MkOPbjJ1BaNSri
fP7CDKZyOVa/Uo77riqdcjrtVUhrm15q19Vbhgp62eXSFSrcQkqz02ArlEX8Kyfq
dDLWlYbKF3bZ+gSsV09fI6FOFoizsJnp5oqM7jbNtfnWAfJmmyrBz4DIM5kDFaWd
TbHpLqvc67nTLEByT+lHip+VR1U7CZKEB3nGME0ovOyuUjWzqT1JmYvmvxyFqH9W
1Cqn9TBuf6XulXt/FdT9TG83SpR/8fxiES0nZI4nOKjC+US6KKhMNkxN9sR7i/OU
NO9PO/+Hmkt9EKaFkTfpLBRXzq6meeQiMRAsXz4zy06esbVj/hxHoYTUamI9RCjZ
UnVT+6/drNc/veCXaSaQO18SSbHemP2kyr/6Vm891ct3MJSZNllQ+gqnkd5E63ZW
HRnTroHT6mYnlYUgsJA4f2sUWkuKnaLJV8UC3u6upQ2XdARfEeO/FDLUzfUfRMOu
OhDw7spd2MJ4rDDFMe7qz480YPzUmzxoNVFbp2V8I40svVCMAiUmtWqDJ5sMu5kv
Oe8nIIVLAWRBEluiCsFVw3CjnLDYdCFA4EVZzh+ME5W4sEUZgWe9hDQv3z2f3c3g
4RJgFpO1sqRse8COYsNZNo5+zPQkiPmnAPzo6mx++Zh0q3qLsgY2Vw4/C4S0fu9Q
NAdC0Ut5VA/F0OAS3ZzQBPXMMTvvteBIkxT5Mu6Z9U4D8PKrNUTMwxalVMoea5iK
Dli5+FsGl/PoLAxEnBbAjLBAuSmRlbApvzgGxE4ecgqscXGUstj/veQ0zuaa4lss
Bt4dm0h+E+fssU5s3Ft2L6AkpzWoprkmuGnxgvKFKRHQWzCtUL9S0qliqGVnOyma
OnqMf6fwbi7JU3oZteTD7x2H6Fq9z1bULxfPbFTT5xNoX3z8n8Q33G+UCtnI3ZMA
5gLNobCmjPeEWbMOduETlNHfdmE4WH7pUuc53uMvlFJVQwn62Odt5byEMViXEOfl
u502JfEQoXIkg3HmfU06sJYK4m3+hgfBY4yrzfqnf9nPxBGSOvG4tj6OyfXP2Rmc
d5Y1f26GFOiZY+798TFK3syDFFzU57DyGNWv8PXavbCOoBqLa4lDEk9xWJ/rfCab
DykiqUo99V1gApBtfNwNM4TDXaUhqbSgzQxcHuQs1MiH7tD7hsw1L6EK4puzMynd
BuajE7cV2B8/j7qr7RQJ+W9YTv2EEU8Z3Bij0BNJckyqHOYRb6Enu4mCxeDC5Jx9
tMtPvo+TRju/yDr51O2FNd2J+1Z97L19E5T1wDRV0F8o+gkiXucTf7gSKCNwGTr4
vHKbYzkW/CSJ3RTAY8QfVkmJb63tzgQ1xVogUevtSJtgZEzCZuJc8gV/UcHGq9YL
elzmGE3WQhuEUHBEU4yJoea/nTat3W+7Ly2zrZPQvt+3cIpnkVa+7YFI5c6R7+S7
CnnOF5rJtj5HtHGxxWhzs9GShjT3z7LXWlZYSWkvkLAhfaQ+nB3F6fgMHiB9yUKS
1b4yJrJs+AbMvflJTq4E7Dge/kNON4nIQEs4goBkSUn/V9VTHuhDk5NMj4N33Q9h
rpVpkm61qVtG/r1i13X443HX7YZo1kDfUonDdw69d8TfA+86FwdKUS70IEp48FJ4
NRgErwTAq3ziKO1hexRt7LKZ5k7oh7ZxNrmrfP2GKMfTxi17rfQWJs8JmRf02B0w
9PU+hQXMKQRbLfff01TIISjt9T9gfcW6nLwnuP5N0d23BQht0dn6kd/Uxbu3espk
0fHHBHtaSJfGYUJ75wfS4SBzxKuguwCSQ4UBUvjieCbSTwgwrkr0afIqh+dCUosk
g1C6OYd/0ny3uiS6lBbuAaeGCM1B8BXWFlkQ+SCp+oftD/kTZFmNyoVL1Kg5+m02
XyBhFPlAcTP81tQE1ygw+/DizEouevC8EBm9sXTWHkb6pW6rGJU+j8sXVBW/j4dy
dOA1BnIAdunR5M7nuJMAA3xbI/5BruWR1zFsDJOVo3iYsellxdAQWBdno6ZvsEy1
7ocNwlwxCvCjal5svV35uJskfgks9qAReYm32ljXmzrs1VRIfYMebSgruPARbbFG
Nn8Hmx/oU3kx4/HWwwoQcY34G+/701HQ9c+2ikSumwbeDfTLLc4PVH2x8VwR6hqg
61tBNNIaQnx4jMtxdkrtXld26hxB2X60QGlBTzbjGVwbkM/hBxK8BCy9R6eEjvkm
iHyZn3qWspSobQC2thFLFz0hfv8L5RestNMiwZc2ZbPQfls7oS0V236KGe2qdekC
A7HLcT95yadl4OtUXkJruASQH5PWNCxPhsOAi8pY1y7PSm0aheMj5P6SurIog1OT
cm64qR50SbDu40R9Ya6bGOfKvB91ctpVVobJAYW1XRo6EXGW58jlQT8qhIOm6YIT
0iMPFrMObfttNy6DrF68KGvXjcBe0XgkPa/s7/2M+tywh0DEc6rFFToVKbeB9bSg
U4twDJDsiSyNjx5/XZZJ/VugKgqACE7K2uoX884Zkttmjh4syhxrUbdCt8EZ8Rv1
SwMIThb/rP3DLAHqgvOowuR8J3PnptlEJ/0mPRwmPrfTZZxjXr9ihiqlY/J8XvmL
9+kf3Ilph1KxM+AExkfcdsXT0dS/PxnNAKjLdBTRv0CAD3oz/hB3BOedu4uU+Lp5
mndy68zVGok568XLEQrdYDRNcFx63lgzKlyZhzZ+IThX85zMebQXFs1DtwTkY14z
tR83wYRDecZEPeyODq2Fr9hKMgrWRU47di3Ha2de2BEgz0Rq4vHJj+1XTjpzB++T
2ZIkR0fWOWwbyqjkQB4jJPjili820lnZthzSuQFGIg2QOo7ZMPS63668fHI8prFK
+zzqXSYwulTZa2XSohoQhe4OgIkvTwxMrRUAwPN1D42Ul4Jrk+jNEF4rhThTxQ8k
mdkZxvfdabeCRToJm9D6y8RyxU3HuznSbdHEdedzl22h+whZdAEqE8WUX3VZqVz0
CLqC8G6XbEMbf51Sb0yMm6Yq75+Kj6VUJMTisFWFKbzwkpLozAaa7gGNAsPY3cSz
ArbTkg+KPR7/8RyYF5wkYaWKj1de1dgz6JjLy0JSwrk+G8gXH7wX/28NAdS7Box+
bL1c1Lge5jIoPbknJQh2Xhn/rAcv0WFpgR8fkx5QN7Tf07b7GDCP6KZFFAKARiuo
iNnDSejQDHWm4W7FWEjTKxHEM5Elk5g/No5r5V+aQJD4d3JyBn7H4mZFwQmwcs/g
v4KzksUmEdjJpHmcdjMFspbpbSX//lUI+i4yUepGo61eIawt30/RSEeFvflN03hG
cObVt9JzUKAcDZI5Z2YTNQ5/S+w6u3mXcR0ShdaUpeHQtp2b9CLMTRNW8WmMYdSG
9XSiY+GNhWPahfblU83A8CcnuA/wktHrGtl9HVcIDoqgCozQ3hTxAoQhab7X7NPW
ijmO/tfI2knTIiDcj3sJmXBqj4HFh+aOfxpbdoQFv3FPqk+BbhX4IXMmLtU+N5KG
pwrJfrTppzrDXQ3qp/auK1Sa4roBg0wUY8cJEyT9aI5oc6iH2/euySoGYcwU0NMJ
lfucJXvfiaroB4VjIqugcefzhpkEuQ4PTikHn7nMZhR03bUbrjYKEbNgeD/HDiNq
pPjtQFhj2vrcdcq5s0FOkk8oqILILsyALK3bjrLqte0JxLJ96QcXuaCv8BlVDI04
QVV3/4Nmo/XsP+rZjub4kOHuu4FPiIfv1n4RPIzc2X6epVjcUnFTFs5HT0kDWYxX
SaBKP2tF8CBtAfM/BgkWzi2qYvH/eoUSfT0LEqVm2fMnUyIXlc+VjsQkk2VzNnEf
ZIh8lN320zB+aO0R2uP9ffY7x/1z3NDLHaWhKiOoZNsrLy/gXv19+qryBs7VZ8qj
nwcBfRD5OQqJbZvo2o7b+F24L8IkxFmKNsHLhEW02y5mmBzRYos8Hi2N9ryK0vQd
DaPB2z+O/mgHVbLgvSobav6xbCbVQmVsguPaN3m5GA4mJti4IyOyESIusorhRWrI
aUzCQeXIpQFQMMmaHqDrbf0yfOhA2kzM5FGQioJlM716QpbzEoJbr0v4EB7lsqvH
36wRkb9GVxad0GSiemLJtO0dQq2eJEa+qbIzGp5gVQMqNP6+cQMKJyuuZWC+X3jh
v92sHd7OrXlE0lCc3DTR0yW9jIqRZ7ug+wwX+OjiSo4vQN5ia0zRAsENlnc7wxAI
6LKlp8rf5INNw2pcP73P00DzhrU7rRBQqFiWfcL/LK7KJu5991gn6dvvZ/+HwKlt
V45ANLXVFOCxS9N9pgdz8q0lXunSUvt9ll4rQ/3wc/rIt5wik7Jeg77MkSXUHLtW
BtD3qLDMEh6Eh/WMIhKkYtpjCnSWG3NvY3L2JD5TggBrliV15dKLYrYcf8thnPQV
C1/AYE24UWDz/nl3RWaDpHSAdiXUcvYVHTqS8h2uHXP7aeEKZdjIKIPscRsTRCzD
15DyNNVF6B8m2dXmKSiCFkOIHadFTQK/rkGPOngn6ZWSOcqNkgqY6VPWQajgvFT0
wMiIRBj2+5doBVoN2n7SZan/Gqkj1UL0UUJzNccdTj797kWGNpnKHzARUeD+bnZt
cx6NlFccV1mUooA/Dt0WZHDLlAbs1N9h4vzLgYomSpQQC33XIxkTRkFYLycRh/BQ
uVfWNGuyhbMHcNTQJT4Br+ZT4wXXwef8/ALnqbF97RYMwS/JAAmsogpt0Xi9r9CX
Q3LLelmwfrASQvcNvQdfMwD7mvyRFCNxXgcngbMaU6n1l1zqFll2DvEDBPZe6wCd
yfD+FF0vdSfKl3GZiTJbXGaOoWUmJWjPHpR+klN2WYXEItwVTWBOTJzIo+sJfrCy
prz5yHnnX6AWKkgIZQ7k1g1wfL8cb85aVBBwC6OyQpsE/RdRf46JtxkAm+lzwcit
aBVyJ6KoGq1jYTSCOIk+9qbd6I5facNScPTKFHaX4mzHJRSxdhB2aWr2VBUYLjPm
XgkWztPjR/9fNbXPQCEGoJn2+zuRqdrSjs6/qvSM0RLYXKW73YS5zgTC+OT5csPq
gVZaogHjbJaius03pw+VbqrUDYf95ir03FpcYDQxRF9JarbqM3AMwvTpsu7tr6jJ
PRowVjnom6QTcfeSriyb8RiLmHjKOvZdcBJyBguz+5IDcWaB8vCdbzwAdUq+k7/Z
s6KJM+QViodC6Xm5Aeix4X68fe0+J+74BPHb/Lw9yPkydKupdyG8WaY3y+QwkN/K
PW6xEe+lUF+1isYKfeoROyV7gnFT9OIzIWqgjsSypb137ZuPQVu044Mnq3GXDgGj
xWKO7enVIz7St6exBQVYFfsjbIB2Zz+1GwszO6Er5HA/HBUfLMbIx98ry1TVqQpy
CL5yyTN/atEc1w9VZlipCZF+8k5oDWeGMTgwzUul9QjXDUnBi9EmGXoPU4KQRjPd
CvJXXhw4nI1hqWu/KIQppa9J3QqX6nW9tubX8T3K4Ky5ENGeVBxgEdwG9VF5wKCs
mjjsqWXhgl9boQQPjdM3EcZjmN5fJ7buDEqjvX60ddtqlTubuOtTMcR5Z5o8Yxj3
f5gH4OzgYCZcmw72rv9zCtwjxyYC/7lxKJ8mQMRe0kGTaknS+TWq1ncLLjKkP7DE
bywZ2xFRr9kix2kBA6r7HgpiD+LR/PIciekChtvgkiUrK9IJHn70qz6jhN2586pb
2V/7oda7DITB41WFcxIFd8RcWhOEBBKFRJDoY7D9CUBx44sDg6yT8+iCJdolIHBI
A85u/TxBdYtJpE1JwRk/hmVBgB76br1+5ZYb/7S6hq1n8IDuCrAK4+hqBsusX3Tw
FAQCX1mwlX99bagz95WyVB6haFck+EGO6vSa7L9mDzrllNVHNJ6wJKX83NSCeB4l
76HzersUuZYPNaj4eV5kRo42nGhu4vq/JuSOMtQvFUwXSVo+chAxZeYHAXJYF1CJ
TQxuBLzvqd+wCpzkujVDyF9tQ/LvVVf75+0djdUo7p33z5P8nvZuM1oZJ6x9p34X
uEJqE7XIhKiQIewU5kpLGluJkhyvjoHmkqyiTV8K6I1qqqSVI/8SpMytlIgdwEsW
GtbnswUkK9V0gpzfMAlpGKCv10KEIXJX0sDJGfslySIozg9BZGrLrHfJmWFjuY/t
rkn2IdiQWVG5bK4mVEbA36pooHkXa+EL6Sen/PZcX6WeGMHrajnGwODIVq14Renq
7xwcj3Qf8jnPUw3dZAtcYN0/JDWMvBaQRU6Rta18sYyxdbRPZQiN0//ONLseoAqM
ld8H/0khjlZTd60N/mlH21eJQuf+KyJbmweflFKGURJ5oZ8arsRQAZZczFqUdCsA
WmNq9c3RGo2gltBdS/woXy+c4HUOx5njld6hBtBzAxK1aBbxyF1RnnPeoYKhRSc5
s0+54mdC91H34hKmn6WH90Q5/1tlFePwKc3LOO+PVkC2SfZaFi35wGhVIsnh57n7
Rb/fS/CGQrbPbYGPNNq0frIlUwOT6QoKsfSssjMxRRJe+YzXuBO3PgfgeiZ5uswT
mpI2YX5q8V9AcxlGXB0vmDSeSbkoU6Msx/eYZuxelqCVYigxvyTV0PljlIDX2cdV
dJYCo0AqWSPo68cs+odA4sn+hAHs/AM55NOUT3/LqeaynkFPnUN9wI6mh+CLLFTi
sKkr2hnC4gPu4W+x3f6B1CaG9dKznyVW2cj8G/P7jQJ5KZOz1zRdcJf3sSTeNmWk
yt7Gr+g1s80FJOuIgRCBLvEdTpnUuUCpvEZXOFE5m5IXFWcIOtFCKD7RwkeJE7RL
5bJNWsTVY35NaxjTZliWypBU3Z+cCNaEdQfDBehEf6BTnvys30gJk6v9qMxcIPqN
ctJGV46TOhnpX9hSZDfU+DJCoYHejIWFOiV2HUBFT72Lbc8xj07ViR6GaUzWUXcM
q4NrAzt586uBDY9BtgCDqKL2tMT3jpmklxWB9Nit1oTzUk5ekmrgvhCP4F9mfZVB
sRTCzW8tQcrSVWcCkKJdni79hu/zSfmsfb3WqRDpezz4jphslRlqtSAbwNJdnAwi
XnF+8MuRVta1hz+/GW1+bIzQX6LKu5wdYKDWC5Ipndqq4EDHquPk9/LNOv8E3Goo
2B8bjBBYksW/5qfcNS78/kYnTobUrdJxS3WYiTBAEJUhaD2AzFsPj30RQsi/sK5h
GGPpAU9zAr+P0IaZKNo3WvF9deUKciPd6rVVsrrRjNAC3GVJ2qYiAwhIUyNhPhP+
ouwzJnTyK1OwfO5RpolktWGyijkmlTH6niaAAjix6N5MtI+OUB0pRWmfNxKkDHd3
mel5knF+zFKdYoLRloXAYZJooeN/v4lEov9QXyIionf8OWXD5TTqjhjcH+Uajfyj
EZTtI6eP/Tc9HMSn9l/VMSuEY0WABwwrCWYELUY985EE0KNttcX0Hx5mITC6AAVU
yvSM86kmd1baipy3OQurGhXT99XHNCcRsLOr+CcdR5PuH9eZBMGpWYr1kH9hktQX
Hv3CoKGrkiCMuRzsYrrqxFbtGzW1UJZ5iJV+d8u3iGiAShbG6JgR6stRCbsqgrs0
CEF9AtwVG1i2xLX3fOQ/F5ACs8pHcMM27L7GBO3gVuPAjg/rUeGZYePIVU9IPHdZ
GN6++bf7gOCIk/fI6zAX6N3haR5CAM50WX7tYgZ769dASZvmoL0IJr4ebWykVw0+
o3HnLcqh+yniu3LjUvNBwdquru/bzbF6enZ5L6/uN+8x7LvwUe0/78HafIEP4gkR
DXZF56oQiCA/EVCX4Kn617hya19h14uF4KdwVkmKTQPhgZpHtrDhgkvjKwd1RLmx
c3KEqrwlwFMYidrTCPrrVe4kGo6AsTRzX09BVAwYBE1Qtw8qJNaUO0nD2NnFGV3p
wk6dMPZpHhXTzBLvtLXf9RHROg3p20culZbcFv+JLOzgzxgHaq8up0jnbFpk1tfW
53L58eI7S97b/35Aw15hHic7eRHiwqGUYSOJaLxlrNioiN3nvGYvp4sX3X3nmiGA
vlzYQhyh5X3QM6D9aKg350XiARni+oJ5zYZZAHzNZIMbw+zcMgwTeuawwPpl5Wh4
Ji7ea08jh98OCQKpVrQuofOlpe2PjuRMiDRqFNCpO8Dd0d10GjPpAbpSLYZjy1sR
NUvNZMi0FfVDQ06mPZUHVCKOdbcRISZtqrHxvHkUjUoOW3vvVYEIe0HaJR+vhCfR
fxfNSQRbJTs8nunZnsl+NhrfbRggI5wfmZU52bSVJGlbM+xcZtm0EHbDn6PwseDm
Nr5244M+h/pyzmApXBxE6L8dGbQIAnLxpBW7/TkV23ez7yHN+vTI42FnxO4HiXAu
B9aWoY/lHMJuOdzUTw6Rr/tX8lTz5MPRmijX3joLTHxirt9sTxMGeieWbiTIc5Qs
rDHVpY+939C5mPltp6t57KVD0scG/7mzR2pRchbt65z5ICz5ljqt2WMkzhLvLir/
9hVREHNANqgdKrC9pn8Ou8UzpRfNDVJrjXQU34+qvWTEOM/W0swTaYuVd1RNgQaQ
AtuWGiGXGIcYRVc5khNuE2v6l/GDACs2Ztu1S+QggOjbs+k8c37nDiWvrBoyrGBt
gPLIXxooFM7702W4qIIMoqY9nbKEqkbZxeDoYcd5QQUg2D9JB06yBpoi7pKdaMSb
cZWu8QYet2IvWiqLsxVFWWDc0dBd2bUo9cuUoLNcZ8nGtowZlo2gugFJd0yCEAnJ
VDEdi6797STYDGJcbeww9t7666m9coiqx8wsfre+ixTGoEZOvLgn1eWBcNEGD3ZK
+jkW1b2jKrxeE8YxRziMV6eauAPfwGaUgkeYE1bApLo5i2YPtMyzs5bsyTMSfLkw
RGxrVL7qLyBWtrEoxEwE4uAScX1FtSSgOCLNn2yUvYakrRnuOE6Aw3pXVHH9YnWg
tFhtnyXEZwaWDXu78c9i9pUS1ksCdYBjzX6K+HcstQJqi03+5/NVo5vRhfvz1/DF
k05LxtIr+L5tynzTVS/7PjJDE/SNshdxUiVMHWS7qVoeh2gA95vJBdOXLQYOxDeI
Q5p3euFpdB540frzsLR6B5yzq2z4Y+zYBB0XnGip+tUEL+ZJxQV3bbseC+Zs+AMz
+a6iz9ZM/EuVAZFrVVdB16yXCb3eerOGY2va/Koavhebgm65UGO/42n5cglbEnEj
WhK0rYAMaf0HjbPy+wpwkR+/e1VF8hpGwxcnsEoZa2XrDkNPWsS7IQWUn/P1bFRr
X/p9hbn5RQ9NATi26IZ+pKVIqNO4vRS31yAY83xApghFYbn4+AD6B8f7QeiFvO0e
yQ0U+ZyQQT0fIt9xGkMvaOySbb9FbYS+i6LyEWlgN0ZQH5Sj1ncdQ7t2a0maLxaf
2xTOu9XAqXS86citMg1Vk9CXm/I6DG7fDejztqyh4voNfuXo6/g2QfvbrxDODv14
vOGvTEXhRBjdBPlJB4AhW+vZi3IomOfEtpjUN4r4Ft6kMBkFT6NwlwFpmwoEaYzz
pI75Kuz2OIjEjD5y3J8V5MWs7ocI3mEr1ZWrwYPOIQg3rYZ+jljO6jtRDI9Iv+Wk
zrvy7/AaL053+5OcZx31rVP+L4t2bGkYifewuvUUkTLQmgAcOG+nzzytqyBzyD8S
Aup1xDDObd8+x9Yfd4zv0yejBWZ6MmBEeyF1U0kAh6jl/ko6WTC6+i0ndKP8riaG
vRxZXnbkxgOCa+f3BfLNpIyt9giLunrI9lFF6vQkazds/J+Bz+Yf/P3YAok+46HT
8bEcRo50iYXiiuxyCaX3GbuSjYxjP5qJs765FQLwo4wM9z2Lg4R66+2++OrF0gt2
jE+N5HeU4MGnM2uME3ALyAb/jgB3RxwHgpuD7I9HpknPXhuA6nEv8vynrXzq2cRr
i4NkM4xwYG4VAbA3l9gSKIfpdeb2GHippQ15L0Wyhtso6KzumwRCCyboH5C4U1Dj
QuX4inwy0eF6qqSp+BoWPIerU1BThjNRJw9ZZVQeT2oKMBUE5wPE2ZfMTwIlv6V3
gDYoVRdyn0Y7vcxGvZ0rMp3rzkNnZoMGWZuRLxcj1Jq9LXGIOhXaZ2vY6DN0I9nL
8zHgrd4WbsooX3hRAdZD6OmnXOIKq1unMrO1yz4lvC6fFrYdvPxVkA+D98oFxFVv
4q+y7Gs6iyx7WgnoFnJS6550hy0Sfd53IrmB9kYSo+McNsb5XVREQznRKvy1ZTx1
00Sh+aScuea3rKO5UaqnItKNKkfJkiz57x1Q4wHuyX1WcNN7uuso+FZDFnrKmkSr
4F8Xl5QXUhS2am7Xs6e6bPO34iD9eg+6998XQ4w8Zhs26fJZTVt+0n7Hr4ZLeR5L
WZdlvEBMnVR0QQlrjusLPKE83rO/oLfUHNTg8Wv5juJdSpdf/blxhUjaRGkO2nBo
0u7vpx0jB39rgitP6r/OOAwNB1rSdAW3NVXmRI7ZWMmCSj4vuyXwq3+yVj8yaEmq
2RuI+m1ivro+OVmU/D+BABSUQzp1YOcRbRpOE9LsvtnhjTwXE4S5vCkYlN4zjDOD
OIftd0lfa3xnQW94SyKoqHwPxMG/wqjyTMAh1Bjm/uUSSKruobM2tLSQxhYDUdVp
xUOvhaM/PR1BukMDRoilYZlliVt5JBzFSEEQitBa9JZsUDUsQ3AcD/GQQxNzLtmT
WW0aRxI8S6mCV/XvpDPhaWEDyTEDMj/0lJed7AdKbJSQgEDQXhlgyD/JIkMYldc2
RbBD4OmoRZFLdAi7f4CgtC0BSTuvSdY/mDUssZoDFn8TC19mYV6YMxEBGoM3Qjvm
qptTWj/870RIXrdthDMVYjPQsakIt/vOeASydWm/dxPAGKaYAQJnov1P74XjmaiH
1q+x8tV56QkZBUIjrEDuHeCPtyL1w3E2S/0+RpEruPYACW3mxnoYL2q7+94rFR5t
vPa2UNHsbiUyghQMdloDRBwzDqC0Iwm/E+gzPsVzQFwBE8xQSQjasSQeAcQLAUSF
OqRoAEYr9Giw0K98FiLvNfIx99YQvHNFqCQO+98d2zPB6BmjoetIZFjX7XsKv7mC
7q/Ir+l7tlZuY7MV9DoDtdtma8KOwJ0UiCKKYw8fm5BLQTJsI+n/V+T3FpluoSbo
4lACdSksB0LDSWB/nVTvj+Ge66hV20Zhs/O1kQthaxA9RfepCYEU/Krio/WK56S5
kCMsNsABPWj4D0IAEmhojF+fJnSm+Qwg8X27MVImSfbpzmRWSfytaGcvQFoD/mw2
RJLkQa+q+FlNx4E0k5pjBGJ/ZMt/GCmOC67wCIsCVKezfgDCOUPGonwbcNY8KOw7
BfGuMB7KUWnSYQPsX5imBQjJWitS6EcGZMrt6wDZn+zKQ8VxZhl7uQf/Mqhqupcz
VPpJ72ahtGjiuKQ531fm9eei+DCx4Iq74Rewxw363SZBsxmZPayg6Qhe1FZ+k7Xo
LeraP6MKrwpEjXtfbF7AyzaQeFweqcyelhp+S0DGaw3/i/GaOa8xisKtXWycHKfa
76lntcgeC0Nf5WLCGZiKI48TRf47fwBs/7UXB/CnW3hI/Bf8D37LE9yIritnMrbM
iTHn0egPl52UeXCsekfr4HHXoX8aY0SF4KNhiwDM88wzqQGr+C16dcbe264UVoLq
m86Hvtk9YfTd4OvLBZyvMLkWrPi/VRZv4ycSSUNufhbTz2yoIB6pchMh0JOuTLTv
I9YAI/5mKTxUIUA4Qs+gFE3ZI5+Rwy7C3mKQ2xM04vVFZWWivq1RYMj4cdetVpxT
fzLWkdP9P38Rg3zYCcz5+TnPXnM8P2/qYUIrp9gpONNnULtEdZVXtkHRzamui5Hk
0yCZW7n2c5tL6NI7DtQox2bZorRIeKEsBCCVc5x6rSoRpLd1K7bCL/A1s87FkF1z
eS58BMg3r3phLw/sD0mXqV0iiNckaDaHDygQLInVybHtmb3RK9YVIPx6a52ETfDB
BwSNkEig5p3RD6YY6A45J7WpTPbtIH6yM4cb5NOgWPzwmWi9afgiZK6jCxYiRMhW
w+uk4qYHCilv6B2sN7qWlTCBg6mWx1HWYH0I3+wHP7fsT034Lm0yney1CDikPWKX
MJNHJd/yCC5AFiT/FKLPcr1lWvPYYwHY9STUOrioJfZzqIh/oZgsywzyS0yMR+um
7p6H4Q/pNXq0xYtzwvyLEKrXcuwb2v9rC8IEBfB79Q8Ye80TpgvJntXARe1AtQxs
l+kzBaTCDmadJvPPYfhRhvnhTdrW5xMOyie1RfrxixJZk9BIBKq8bO7hAgfIx+4h
RZu7mdzZ6IYwXEQ2mVw0PRcnu+mRReCHtCIzTSINwOuHrABbRp4oxnJ0gTB1xyH7
keyIMlkLu9MsJRYvlyGfEifsr1ZYnTwlZ3RqkYQucGYmn87+sz3BdniDsDStbpaM
OaBPkzTn8HH/3kHOeEE8P4lx7bha30rPP0tJXb++plk3vq59216jLDp+8c5R4Pfe
NMbtCeZHbJQ21fDdX1KQ74uWVA+M3l5+9AhLR3qevRop/ZMxZyAY6lWQt60d78nk
G40WibwRZyE3BNxKkfcAdH0GbN6xNHThICzGFZ8Q+pQ1C8yBiVv8wp/K9zwUwb1R
s9MvH0Aicephf0FTfhjPsnsSmza5qw1tagf3T5NPwXGybjBHT/WEzz0APr6lZ4mf
OPUwSxvSARaOFxesy3qOeYK3VxAEkeRrBObqA1f40oW/KGF8IzU7HWpupfMduEdc
8ILnEj7doxobXG12o2bsSEzCs7mdGmjWBQGoribOqsNgzPBtLG+epScu+zA6GRyG
0t0tcYa0VEOusyXCjxK0n8X8zh6Z3D2FLQkBC7CoZK8gO/m5ZNoARNXLFzAmiKtl
spZfihJTRAC6mwmkvpPqGP089LyhG/aXaqPMw6UTibSNb++CbU9FJ9JWNmTP3nrs
yZrCR3Lk2LzmQtLDc5Ctebsqfn12UFwuWKklUtZm2l1+uurY6YMSG+nqY7sW3l77
/6qyZ9WRNhFwW3kv/Cic1+bY93wKuwtLgvaMMDgjDgrXU/UVZqczoNzV9OpFirIJ
OcYWET4as01StvCvRYki/3apZJ/9zCLs544zznPBcfZV5h3R6ar8Dkao+ZcltRy8
Vc1alRue+OLpHISCfah/8/QYPkLbgExScBtcOrbHeZR6yGymgBErzck2uNXyG39X
usu0z3W2rl/YL0d48cGHPQGWPnQ4he3/SOUTcuRkEQ1+g+qywPqwZPKtvWpAnlUn
6nGZGlfY+rHqyeFaBq3KPb2wq3Cz3ztKuB2/WJJLvxwvSg87kBnz3+VyZviPJuNA
hOMghBRLZwAPPb8uxzIX+DZb8Pe3E1/pswFfzCOiXdBMAs7c+J5nVDmgq3EzUuOr
KH8CLHVUjXQ+TtOAKH09gjgBxnVQUcXvOZ5mSBHJcyhDGHRf15eHBR8Pb19yth3v
kbCk4XiEfHOQ4eKQMu1zW4dZQFrTv63Gc0w6HsPIL3KGp7iWjJlMT5Y7nldj/JSu
rJk4rO9rRhJ26nKKXmzVYo3Wg8heobfKXUh5/r7+h1DoRDSPx4wmYHXQHWcMdHC4
fALdxQdbi/10rk6NNu+y34WsACbV7vNBbSJ2M48VXHw3pyLG12G6u3oMnaZpTmdG
E+7trZbC/f+SnQVtN4btx72p/9/MnyEc2iWMv+Bd5To6RzphTfFIJhbrMpuX/2D7
2L2KrdyPRAS8RMepqxvEaV1XHPd419Futj7BlJic1qpV6Q4bIjQkG/PUhEWMOImE
UeQ92ICi0s/H80pWDtMCXZOo02XqnlHbY62PBAndU8X4MfIfzd/zCn1fqVNwwXXl
BPcSNwXRxmGIkPQaOgmyqA83XwP2Dwst5YIbkj58Hb7psFI9vj8wckXah2Jgrhlv
Hqh6FyjW8EZcCSPIsxxlYOaGV9fbCg6S82Q4xuxM5g3X+P6ydnu79U/HMz6Rxqhi
4G4TFwfqNTZWQnTjPrBf9DuZbx2KMAnTf7F+QFNEN3LrIYMj3pOLHA40Xjzp5tg1
XsFeYNhh7SLnSgpLExq1pQbsRV4W1OPNv0lYzDLn9I4TxuslHoujs+2vRKZgYmBr
pCySn5nx8+wOqFOzrzYzOVb4oDpyXCpb2SF0vWiNonaD2thD+ICp5K+FCE90n0ip
WSoFQY6JESIQgflW2/2IJ1geUUBXVCFa5C/+9or9qXHDPCjQi7VVRn2PGKLOzGAM
eA2VATOafjVybqdcGiJf2/YcPqwHRU1PWI48zqEZiKsOlGdo3VXnuYaFqsVEIe8X
3rXhBlYaHb6QK+iya0q2ZJOl7vHhmdXwQ/z2Ui4W7gAsP5wxjTlQ5IuQhx7oPHOe
yHfaAVc4yVOWtk4hIX9JDF8Ul9dxBg1lWqC+Gf3kvXClefFRNcWD/LWc9M4TIzIl
47BLNHVqyvJngMG93Kq3DF8e+90Gpm/LrnRmvNK1ZWK3x9jQIwL9ILTLQ+zJOzpM
+Z2iMkPK8ZAJNXSGaT1iHe8fPfIyQrdfnnu1KKJHFRPtpqCs56B0csJxHq+yAsFC
u+Ab3ldJxwcAOIe4p9Hef3SE2lhT4TeEDVuIHcU3q0fUJ+fddCvs9osU/DDzE5tc
vwdEG320Ax9cHBmCcBLTYxDIVDIzqkQnuvywQLaPiBeCSkqRuEZpjE2JFasKYtA2
nKi1SI33ee/pfDz4cHpbPimANVE+YDszxTPmSbNMfW1aOllzlM37D6h5o7S+BNCT
HYx35JE5iQImy5ySTBWdJ7wxHdVmHg0zdggkDKdtlUg73dwsr7hLFTtcDex5u19w
DdrKQ9XUPkIdrNTTA/DOuJVwGlhNrWr+YZIBslk4v8A3jSSVsIgWOV+UE7wzLPTN
QUxskzfpQIwDU7eVoPsErHk/xKWVanKoQ6I8HdGxBWjkz4b+pUOuFNvhyqgStYud
LJ1bZGaEV8BuKOZmAz4hP+9OisVTUQzDi2YdtJeTKozJPyd0HBZauypIjurIHotj
NOgoD5CEWjMeVA2HtXoInM7ClGytMgrpBI7NVQx/un93FtXamKGyfboQTG/sBpUi
tb11XbdDgrawQtdhWXb43UHff0wc+FJIEliz9TinG1e4KmeJ4BopFm0OuLWNoisC
DDgI1ae78x7QdxTkwgVLHDornheY3+1sPoLd2Wv7t5jdeKo4+P/7TNr5TL1m2TYd
QLAsTaY0ICxy5MKUOPeC6IzKyGfuQWCUuESKLsY0/O0i00Qbpd0UjQ6j4tymII2U
V+ORYnxRicS29TbULu1Qf/yasKyVzTGYHTexbKZcYmYmy0/2fou/V0Aj7D4JBPEf
gIrWfN0oi0hP5e8MuPou9G30OGqudHpedp4SpRoFeNGicjAA3+/O7rearZI2fEeU
iiAPsSHZ8w10JkXf+kZpAFKmUAzDMddy703oVoJxbauJRtyzVSyvmde0irehdFCY
yetmggxwUMA8oe2tFkuy+UY7M1ecKAhsQ2M0yb/elzE78s6A3OZP3ZfDHaFFs/A0
VId0BxOfHe+qWdr6vopypdpuBW7kHJsYsYgSyuleHPLI9UUFh8LZDf6IQ92nHYrR
GmfHJ8TM3DkBtcewMSaov78UjCfcGTITp1+z1+dWHFEjBd2aBSwdwJ110+SNXTGG
Nt8k5u0kFQ0a6hS1z7/DUiRSHt1lH2RIbb25o4PX1MqvgqVHGThlP86AZKJytzSW
WE0+EvCtcJ1G+kxSZX6JCB9zlowrcGkoPNhqA6xVUjRFOokQ668ELgtR5gjpx+dX
y7l9PWzCcDvu7AmkL3FrYnvn5CW797rLlE9Wz3cgMFYrPb522breiOnJa5ZbtW6L
FuFu67ArYF44oWTsSXBxg9u8WnSp7Gir1fLiviEJrgmIkmZHDc499K7Zw/SuqDPn
t8G1oxCEVDj0uGgZLOiK35/DOadWcd/wblVvd3Te8Nt+3YuCDikjl8SyR2mRCHQT
CxaR6snLFc7+ofxU6PyD5qLqd3Bxop5EvYcuq3ApbKHN9OYLqZAnBs/ehCiVaM50
HFGAOqjs8os5LJv0W76tW3VSggbuys+xdPQ5IQeWGQatOC1Bi7MyZYh1jO9CyJ3Z
p0JkLMnKijWhE/PG1UhJs+4e/1Gk395LBS1GbxMIidSsf0+3OIWh+DOi1wak3jsc
pFXO+w7FEHuauvlvE3Gvg/rj0i1qxxF5t89o1HQ8ZmyLhcKqjUX7p6ZZttz2BrHm
XdTJO/jTBvvkcbm0UWFp34sLwA+Emc2+rmnYZA6E5ckTyhVaRsg8ss0jCmf8HJyS
Vq01GJRYDNCJfsCCCI5XFinRipXpRPUvbISYh2G4tkrwbkR8MSMVWM3TDA7yEs1Y
Wbyn9bNydMgyVfOjSniHfVq9URBGBKzo9zq5kS5A5iYS3/fDFVG3GmFRKMwfgSrN
vs1qvJm4hNSQT59Vw0cM4uoC6TVwGLeAwRCn8BjRPXtx8hE4jNCj0IjdeX+5git5
ZvEG5Xdm9kACwbpWlcLKsONVJqcfeyfOPFthEe5PypK6knvHtZ8vAOdoqciPRIL1
G0IHRJfuFzYI1BDpL8qH6yb3I6oTIRwWDdCewuqAPCypk+2TL5TFQc3Lh2qeOjue
L1YlYL4ULSfA6CRJXsdt4Z/LQ4emslBDw7ZABL8fOy6zUPpWtAmcw4rmtbOsxEug
uG7BJlMf9uiF/Iz4dXPDZQ2mIrpO7NE+iT3sSBBK4G9IngI3LEYoMCi/DYm35CeK
Oi8Dyj7fSC3k4ZpUyKAXWUP5CAcbwjwAwT9yG+W7zZE+18mD4v+TETn2T+LCJFrW
YGGPb4wNtlmeyH2gkH56x7tQKJNWJ8Anu/BGaFhbcaeD8ydFcd5u99XhPHB9d94Z
VtThvfltTVPH3vkhNShslmZf7dCH/L+8+EqZR12QhilvP51jFq1Ra1udKvefmbd5
W2TPUl7U1w/Gi5QEDY/EOQkAhxaBqy7198hfBeLra1zL+0FLjfaXZamb7gpje01n
Z261nYtJ0Aer4NcuCDNKAHhjzMBOjWqCEuT9J+q5M6QB1+evA5goa7TBpr6LXXKH
d5JPrt0wB1M1YRmkC3zJpID5Bb9f4TWOW50JukYU9Jv1HO1/c1CHHZN/zk+3usmW
qtl4VURSl+dZavO99OwE3pC5/MGFl4kvQNtljUHEWknRJPNrzRpZWIH843s32GX9
03ASeuVAdhq6nBEWoyQcslSvIBg3khT8FgtQv9nkele6iGMa4IDj1ddeUPWDJxcZ
aQxqCQW1UVN7dsTovCbBxs2jqQ+19RCpgPX6xD0IQZ53PjsvT1CbLo3D46Pjs303
5GZYO7A/00nIh0cdZu5ZmmhfEcJh0H/ShAxCnJPHvjWEA9DGOLjSCYOe5dH1BtOz
8JRlztj48fxJm5C/13CwnNAjdSm+8CQRmiB+2ZNNSLDClz3vhgLDOAdec6B/AvBa
QsFenwsu0gTHSnxQ0SiM3pPeeZFjlcPzDqcVpa/gonOlDVVBBqNtem7QTqMUJpho
gGKiPRc62nNLKU0pB2Ll50AvpXO9C+gCaGaigM+lf2YPi2LMZ6bolynZm34dakIn
tvmJys/FxOgOehavxWv5dG2nCZ1GhfvdaJI1EXlsfAdb+UDvqwwoYy5BL0ngoiAu
uxHOOFztX9HD4fBPKJGYcBjOrWXMKwEycEoe4vd6ip6TG/wHyGwwWEOwm4fMLM/F
aMcXANlCy460AA5WOCSJPwl4lhbuwprs3WnDqc/fJoYj7FEvJBoQhgHRQ1XuP0V6
Ui8oZRa9GmxqlHEST5U5YN/Un/C+RZ5+Ut9OPSk+hxFluDhbNSMtVY1h7UHvbDy4
rwwECmJUKu1v7XVxLXc3R7Kdz6TU7mWg8u4ZS8r+gaWkJeKX0XFWbj0Fmtr7jQ+/
xjQxRyx9NHoVAuVZTNRLdL3RFbEJ5F1l6vHu1NQkG8Aw3Vff7lX4a+R3ORbHs/mI
8IGgc7lCM8n7/ORbejg80WiafHGRGtWvZupaJPgHAJIN4/HMEJx4XaqkOrJiO2i0
9fUghTOYt8xhdAZbz3zuqBG13syC/7uI4CEez4LgxM11ias4KmBpt4wZHyEpY10i
d5ouwoXdrnPyvg2u5nFVxki8DqcserLwjYPj41e3PGE6kSxvTMqr0Efqc8YT0UC+
43XUK8GPuTy6t3saZ7KW4t5pfVUZ4qJAd3nTCJxgEM5UgAm5pcb/VeMMh4+5CyJ9
PCUANpRojQpFDHrYtWVjUBlDS5JuQKrqTOeGtMXcbSrcTm/ldHwpylySSYizKjVi
LI3relhtnBA/6j7faIdZAp9dd/d9WG5Vrb6OkypzlhD9GjBJWaYeLXdKjiXWGx05
wsrGuakxXe+LHUdHDnJ1kDq4YxRP3FRYCA3GE2ynB+wn6xUH5cOgRFupNS7BJORf
GLz01E6P3LB3mg6oCXGAYILd/Wckey6Dj10qjAWWOlmhJ7H1DRNJjYmT03o5QN0b
iwQQIp44dVkW+IDmmDeJOkXPFS/EjKLqnGaWCddgeiW/J9OE3th75FNSMAJLTjkw
WNg0tzt2+eAVPqw8O2kXRrq3NyiOMcmG8y/wtE3YbBxwL4Rx4Woa5QRVcRBoLr/M
3LzCTKUSG2VUPSGlXVNoQkdr6gY6vGqRMYnVdt0CIGgg6C6AOXM8FtQD59QyMGw3
QemnPHet8Qz+Aq4Jb4JGT6SDVodnLBOYPKCw6lwkeEdEgtwkKeNbKyo22fUkwESb
D6K8SldwNVeeMU/4ZJbKXie5Xpkc49twP0cr6bzwV1g4J33v39dyGn3YhCvvsXQL
J7ooLgsGMlgmuKobYq1XMcT0q05G4DYv7L8I6Ghs2b5ucWp2MIg6zUVVLyvU9jeR
L4AzKitjqVB/mgKi0xfvF8mwK7aZL1VRmv6jLLQ17/TMIvFQ1ukMoVxl7Po/rGXB
naXp38mX7Z4pWC0yVCa5HkIt8TZhtip0rva7tMsVbVlgx6k+2JI1yM63AlEWT/r9
8AAoL2cvwLo0JomLmGineC5NBJnoU6NksI0zuHr3SDXUmI4ImEqtaLEhzgZSYI+r
gwne/f1pe3GyYu7s87r42yoo8cRwrFswY8/IYvbC7Eg+HGmSp/7jP5TZ985J2giR
7o2VGsYp41FFxyJJtRSA7wlSMTQQETSLaGWtozu1bOuDofFeKMOG6qxA+nim55n4
YjGKJ1psg5NrXFwURvqg2cN0wtz0vPLmSwDb8Zc0rklc6TuSo8ExMNojUqlp/fjg
JF+cvtwJYFczlWXbdIb0eZ7wzKFnk+PTshZQEI8mcDxGSoLcy9uEfO6ix18Gi9lE
PejVvQAoahMZNyOpgWJRMcX/W0sQhxmjsf6KzMjetE5FZNQlH+ntE9zvsoqV8DmB
QpI7ZpERjV5Zw/TxKzKokZcpddY60/hxXaeZHWX4PlHLW+WpxbaIY7zcbJumidWo
yD5c1i0rOC9JgOFbeGeYI3L3A/LKUQiq0o3vIeOWOL/JL++zJ52jnrVA6dPMqoiL
y5W+sJOAc+GJIpdXWfaUFINLjPOvGiHCb6Fw5HgIPrY18AqyCxeXF459RIwwjTM9
uq1JF3GEKzbk1zzDVJHw68J3EoUeT1jdpnJktvRSGo/SCPlgxHgqhL2VnwxHpISW
zM4wyAwWYx+ooajR6jbsWSYopNt+KRAiseiqstxlfDMuWXav9Sj0uumH3mpXw1s0
9nsd8vSXyh6e7X4dT9trK8q5cu0C50rQ44Oa97UPIaGIYCuvz2W7OcI79sIFGqtf
6+0iLhMz9tNgdMwlspqZUakemy9fGIDZ3l/0YvdC/k29AWdLTL00NgKePHs9/PWi
qesGAUd6Be/ATzAFk0eMPJ36YYvL48YrrFbhhLQS4+GK4Hy2yKJ9H1zVBQBXK6Of
5UCnTxeICgITPelCuMRZ2F/8stANrkXrve+BX/KzlWKQp57QpO5xpL6v9GK/OiO1
hraerLOOYuBJmB6lVE8i3E41E4dtEMpWu9iMryVy1YuZHcXj0ZEbk+/UQwFbYWyX
0c8r+j2gjf4SsyArmcuCyPQBOHT87TTL8JT9JiFVHkyISVAB6Kw2ZYoKEqvDFtqY
QPSWSHm7Yl+jd66R4jPJlj8e4trAMmjS9KyH/boe44opUMQ3dHjCtiraSIhMhyqi
4xZscVfsqNQS2DJLM8NSRrTpoxl5J9vyEyCErNmTHDZrKDrHIprs9EM+bMWQVme5
4aX1hkojeMkVEpZ3M6BdtCx4RtY6jjM8yI3BON+bfP+z0lKffftR05ZWtnr+oKxC
OKpqtm0e3JzZB1hDby9v8g4xvBAv+RzAPMeR/A3MJEeMTr9UKyyRkyS+CRNELuX+
JJIPQZ4UJAEhHBsWy53is6hhRHZ3+euQUXDpLTvzj3xjzbJ5M812ZLsqivttMjI3
G4rpdM8hXs+oYCfh5fQW+gXkQ/O88AbjaMvea8LfCsXIMvVCSDCl1pJtiYVTKMiy
2o/sDw00mcjeUZD/oQApSkA7m9+RICDyAhPx9Sju68QhSay8uBpaxEeCmrMPDZKm
a0CxqDkjOuX6L/gc6dQB+qQ8eWcSlZ1dQ35JxNOGlS2EUQIkG1jgeM28jEtUeSep
4VZNdTkzFuiTbYe87+he+J6wx3KSfGOVv+GKE8fJO7/FF7LvsqiSI+K6V4aWlwoR
WuWdiI26p+9Qvu9lfhndTQkWnzOyB62HUtMroh6g5nQPAo79GgkqkDOYSORD7jaH
cmDXlO32EHTkQJw4lhHI59juMKIPKvSphEKEYarxm8oTTMBAOs9M8YUyZB2g4aba
3KOLf582mAct+0IWWPQMCWqBTPlA4qs8TWd5KlV9IdbWOxG5VJZQAZUyhQ9nrs5D
uL0JNaNp2HLG7Pm/HWJnfjNAag6qYtA/MWNqjwpqGZsaw2drUQF4UiH3+RIszIlF
/iGQQ0Y/BSnXQvO1whJ4TWvQ84AxlGkbTSto+QpfGniLEdfPFUGPqFunWiPh0WlD
HodnUb2cXJXb0DEGEWJbqeKR62GSZdokLg1Wca3+igDWDwPBrvPbCY3bBwfVmjnM
Fp7RnaWlhX6LFpIfz92+/pm/FGC2B2zLYQJWxf/slpX9n4DEX3m9Z0rH5DdQcMh3
kcXH4FevS2Q2ihTI2MLrty9V/VtpqIsF+Dom0NinR+zAMdrBn53WL19OGwUelGCE
HvtbhozzoKdf2qiqts587KGsItLIOO5jSZhhI7hx5ar1lyOufYCd87+dE7+cVHtv
u4pPW0BcGMGPsm9jz/g+NM+Kb6RUECZIrxVgYLP9bsnFPyDRumSns5ak5Qmo19GI
pOCDzy3N8GFq5k3j5hBkXE0NlJAMKTSZfoZYqQw7cEiUr+2fAHyWtYc1MA2/Bm4s
Yuws21KPWiBIYH+ivr0ENecAFMVih0tYPZ9MJpRuuWSCGlsncXuQ39cEU58eNWXm
EoC7QmsLe4UMigolZk0i8zdZdNSuFf95gf9ftD7m/5TQM1+YovJtocQ/IR1uwAVh
3peltIzTHRA2xEvj2iy35AQh1BmguiLusg/p4FMF+0ubcoM/zeHqpUVeOln0x2du
3EgVcLf3wJMCgWaGMtAMuQ1VlY3TVndwzPRKH53+cp3RID3Av3jeAeQDV9WfILXB
hKx5PbPaAb1LbnO+1Sp/B4JNPIoDdmAQAzvovFPs7uNAG4qnWyUK9uVtvKXqzcjG
8OPCIVFz5sdAsoZW1hcIYYiyCObJWXtTLu4vGCgStY05EDeQ2x5Mxv/1i7tASSoL
7QwbpZD1HdvZjTTr9tAlfqUfmIgYFjuN7+9fXOEvnQMWkDyhhoPB30SZu4S/zRCM
jdi5AAiuEOYSN0SXcPvVP7aLatQAaUwnU4QecNyPNxnUaX5Dg++h1kJGbY3xmuYz
3sO4CxQxEnrQWqnAMxQDVVbODBERzTivck7HVkt9CS4hkEQrffy3A4YfWDoknEgH
5eD6lF4q9z+PCmR0HZSsWzAgqFAcZphC+9sziZ3VE2QF9pkuR/zgRlPH1AYy/nQL
h7pHDvbm+NDji3wQErvVl+mYUf76ucZr7yTj8seOAvsrOKue+YfJJbajRLKunS5P
Ro3mdfBatO6lYWtnFllKLyyBYKrAApKd4bmowdOuEAGyQ4sxEYwlNkqNb0KcnGv6
DLUkk9L9H+JIetcuDCeklz89hJnI3+64vMekAl618ubGluKvS1bSLXXveNBxKyti
e0mAHdZkslnvlfwfNQmq8xqwSs3L5SF0NwAuPLVO9ZabdDi1AiQ53ETs4X6F9K82
4Wmsk+tG7+BftO+NHjlo+ATwCr2ihbmnLgcPalw88BNszU8t3TxRbBtRRpa2OZTU
1cqO/2xLLehqcO+vWVyf6JdX/vle0wpZlT020dvLgmhayx2pST03xe22ifypNgJW
RPfWWUWRqmlOcv3G5DiB19yum0SJDMjJC+kYeCXTI16hTRD6HkAKnY9v8+pIQ9eV
3FWM7LN70HGgjoWeMBuMkLURrG1jI4pSgytaw22uYM8BOsSxPJoy4dtHTgxqcKI5
6ujLu+4nBnGVc1F8Dq5Hih1TgvW8Ikjja3mn1MfHxB/pVxWa7Ag9jhtP8Eq5Tr+P
XHCPGJPmtST4bes1/iJkKRr4BhoKQkFQrth9L6nwvt5RdRoS5cFPOMV22ZQXfhvh
iHMTgj45g1yDK2O+94GYM/abHhQdJh/lTiLlc3p7FIj7qXHE1Wq5QDU7dC/GciJ2
Te706mTuDZHjOCoXItpZMVT2EAbLckqnd8vPVvkjOZIvEesqGoeW1D7zzPSnIFSf
gfdkLvP2MN69V7zDEOQ2CrOVxNxiYwjbUqE/3x9y1npKseoiMQ13Y7C7bDFB3nwU
YIjSDEf4+VfwYbovyKGiCz1z5mqRXo+DkOyh+dN2BKpPpADWZiWkpz5iaxLFekE6
IEGUvCyC/17apywQ/PanuzVMG2IpiVu8EsoKv9f9e59SILZ4JArX3eR2ENtmEuNj
civqbLtXhLtTwsVxtTa1CetbppZ9JoEytr8Y1QA9JoDAbRfIRCPUqa/LL+IKJY5b
kjyXuRULtTWFnkn2IT6YOLTBHz9f6gzp69HqRoWDtRViJYxsZfnWDhLFTJ+kACRv
t3DwQGBOTcyRm7PNkvFfvjPO5IieN4PLWPaK/wEMDWd6P6itSNVcTX1m4bAvwu7Z
6FrX9fEXD7oSNa+M3lljKEVTg0cZiox9+qwYDHhqoKM7fe9HBK6qW9KTDLJ+9Nko
PdtAlr1JYCzL6wiTCp0jdg+fGXzmGANby2B9A17lhIxescc1m85t9WRk9CTc/aDk
lzopZkeLfeYtxzH1g+bfao+UwETUzkCkO537RcPxj8YrRQKhQavyXHxi+kOAbdcV
f2xtV78xD+nQmKXCgqerjmZwNLQHrqvJkFVZY5Y2M0Xk2Bl/pgl+KDFH6NlhC2GS
bfMUG2Pa3+jh0820ZnD0PGNVkgidgodHoK0OjHq2CClZQUouIb+ZwdKWzvnNV9SZ
zEYb9PS9jvKvR6pVcw1PK42LdxWRKNt2WJRcwfdKkbhtWh488tG7YGDXXwr0IJD+
i/n41YxpGwBdNFfGwufSOpn6viHbaJRxag7oa05x31xubnf3b/3X6oVXRuoSboI8
roqBcdgugLcKd8c1rCxnduGtpyO4/pzVQr0X9A+lPi2jzmmoUC/iAdR0cjz1bOoM
IM8tzuIMNIG90vpHBB/5kW6GjPybm3fs9RNvlds9U3QPKsd+3OdvS9fy6jA1GpTC
CsJfoC6bpdiwwl9mPPtUra4urAmZ+//U+m2bhZq25aZTJL4qn7w5swgAnJnrSWln
OIyBaG1h7tX6XHILPQvlzJjRkcwZjR8ZSzgsPEb7bKul5uW4MmMcxjdJWZmfGl8U
7kclomXpU83zw79QqzmCwgr6z4+5MO/ben4hh8WQ8Cp783IaZfWaBsy9COnB+7SU
Qc+F9HDej73xLccuL7imLNeCrHCXvOxM60jPeQpyD6zQW0Q8A7lq1cOxMO7VvIaz
V+WtyFYc6L6tuBP6uxBPT+/NEWoYZsyMo3bqrA3emM0XkzNzvErr09/dU2QAj8Wo
sltQvNBSnkJId9kc1g/8g0ATk9PD61T9coXlXwqoQI6ymDZbvrCMDW32bgDTToTf
+1VIMcnct0ivp4WbX5McOYNbzDsQZh+rmrzJ9abQhFfM7+fzyQxzARakYmvGrGXq
ko5clwTVOUEJJoX9TRuod1e/OwgLE0Ai6pMBwK0gV55t8S/ppsvcduNBAn/yPzsw
S8kMmEDd1xPO1J/qHHiTs4oGifsK003EayfR+tDrKQBDoCWLHdupGni738g7uGOU
Pc4wH/2NOoR7vAqpbi521isv0TdpoSOmh1BivRDg/4mL0U16quQjBvKyoYdEDQxQ
h4bP8vMt1wYu/lxWaRRwj7Xa04yqKip74BHHT3jXXZxvd1UlVrX6ena2GZW51HIF
j7ONflCtTXmmyvcd5JSE1SuyWZMDefX4K79uEmioTXoayhcMx1MMI5b/rlV5py4r
3dqfpLsByXO6qomPZRQLWPfRVCrZ5N2S6KqrI75/rfWQhu8UWhnxf0rGbA1BoYgC
XVVjB4ioq+Qa/+afyu9LcBtdsxF1rReTzkA5Z7/pkxvTQjYIt11hrsZf5v+FBTMJ
ACobRbO5s8zkZk9AA1yeZ4s6DPVkbS5kT61GorJ3VW2unP/4Mc38o6yKtZKaFZQI
e1Hbl1ggptH+yZyiS1lTv8AbNQZstwYhxs99mta0NCYNscvYTd6+aIANmQ9yz1XX
1C7G4zzGlW5ABKV+yHTJsgkMJW/xigqYlwxlPqyJlrsTLkai/11DCd93ESycz7rz
/XC8OnEAnrNqMXm8bqg1Bv01glkdO/BpUOHg5KU4rNMmX6wXs7a6nM622aaH3HGV
xZNTzJBZfmXx5N2RZhAYJ/S6TOzeXttQF/XdH51nu37usLBxF4UvDkZ12C36E/ym
pWf3Unrl/T4OfDp+YZneK2DjjonAXjC8YTDweejyv9KaAnN63j+Ktw2wPMXOVvjQ
UseA5QshuT7QxINVJis9d4362dJ653p+84jG0YzLZ2KyCicxCvyVAliGQFhMG93A
rb9UXsm4Vx0OIjWEfCKA4Ws9bIM9/3ZHD18sbXkPq4hOy7oXEOTRo4YgjT3uj54F
G3r5yrytMYNzmVmfnhpV/enF9oFocUa4xTCrGCrKh98O4ZL9I3HTvJZ/m3JS5cyQ
zJ3+y77tm6XTIvcWri92JFc7l2A5pQ0mRXlc83d+vWt5mwS0mIgogxOAMVLyBYCT
ApWxquzwxFF+qb4Mqrdf9wi09vPybi7hJkHJXwBkqWsrGnyHkbmYDCWhmrp7mae1
yZtTyRbrt1A7KfZaPvApPm8GgG05cO5WglucTgBdyrld7OAZiArE64/vfT8B4npx
ofYDAcF+LsmAnpjZlAHNZpMNKATTSsQX9hkLfcySTCAF/ve2pluehWQp0SuTqB7A
4UM/Gei9M41duI+lYshLpKHOkPjEogSj/PZr14hKlYH0wup3RgciyDMkijyKJUAs
RdL0Il4T/gNQAI3Hsp9OBudc3U9oyuvHrsl3jt2k9cECh++C0IzUgp84LYFxb/tN
sWomGASFIctkOZTxa4KfS0cvxexCfNv5z8YUbzE7OXflxrXVryDa3ajc0D3IOyun
z6jVhAGqD2cTjlAeaujeMLPPUg+mcp3PTtuRa5KsteBOP7XtNlTAtiNNsKlCZ4g8
4TzWdjnPyGteeSs7ikaTe2YRd+pgyw0JOXdbKd5rF2wLFd1fZFbr11oLXeeWPNM2
G7pLosI0LxeF5mBwYtcFH/lUJUS79VwuOyx5JWKVRi15GbF/28wiKBJmFV9arP14
BJoGu66FuUsybCMDQwqoylk/zMJ2jJmy47c3kmGrG9rmLeDT9RezI5PYvxKEdVPR
qtdUGAVL1EvyUZYmfOHuQxVh4qnAMiqDqEOHOOrw/1fcsrApGOZbz0lbYqfTRaKF
DFeoqZu3Gbvm+b6IVRvuAuXH/LnmkA1r02TnDj40V7RxBeXI9h8AfdmhY6vBwV5i
mvfyNDpceGaJugUJfbZW1PYreodIL0pw1qoGHg3qh7gKigG8SqLtirznMsfDJ8ou
EB9b6/ccyuLIk5vr5kbOZyLa6DUUAneNbfgy/7h1hLKE7VgScK+E+THUbmT71BSb
hrOYylh55GXb/kKhBQBy62nsrqsGE0mOsmTgUChu0qZKesxGFCU741JubrLREh/Y
jwhTBQhF5IZ58iwRim4MtYCSFpV7hXaTpIzcJH5IIvsAIyuKHvQLxi4ohaIfGEvX
L932LIV70Co/MB3a4If7y5l31AfI1BSDmKs2j2W9TqUS5I/HfyoFN+knvx/GzsoR
UEQGZIHAOXXficM2QrAS5hr4rVJUVbZGsPrCNUg+d4I0j+NlNuCE6Ib96mdLDGEm
EsJWFKY41T6t2zFhj1r8BQhK+kQcSYNF3/IazveSoNPsZQ+xI3DRetTm4nMSW9DV
n0HBcTsqVl9E+koe8f2r7V/9DS+XNRVDUdtFAM5tNgqUCjgPnIM/5JkmuWm870WY
BtRCI5n4At4+m5jhzgHVoVFYOccXYd+h27UMw7/y1PxQbm5WJ2+DU036BrBbHcu+
9gG0inar7Q0F6oGPN7OFULJdCIb/BJ+41NvOxGK8k1dGhYSVT1coXmkjPeCs3O4m
oQiJQJJk+7vAVQPjgrntTCZTb01rA8wban28RTYhrGd8fL475D/4NWO/av6Q2wCF
fwnGgBesceOEIvCBvVHo3EG6L/3vS0yOKhrTq6ohgEqhaRMoeRW+D9jSQSTLZRGl
2dAR9eY8NFckINNGHkmd72yABTCB537dcyxzMq2Gz5NMbbLspkgruzhUTOIV8ETk
tksyf4VOmjIpyCyfnYdwKJtOkAqLSICKeliqE4CIIDsqts+PAnRhsSI1WtxfIezz
aXknuM6g1CGvZxqS1cQrRIFoXjP7ZioAvFSeA0Q1FmchyQyDm9acfGqAr+K754u8
U0xlVTzQa323+OGxdtnYkFa8K2nrc/wyWBZX4cb6LlklJDhrqk78yFOSsgMK1dQI
i4zVDhVO6DHYsjA8g95bmPpcNmH1fTH6sPCsRsnfVvKLhkREKB3LreBT4t1l/3ju
vLTleWLVemDWwo0E8em2VnP2jLqbuB0KMgn0ve/UzJ+rENiY+K7lz29SIP7M+EJ/
VS7gFwGQHhX5oCnQ3jfwOb1y0F+EO5U4aP90cFdu69spn6ei8oNEwUwm9+MveMkH
c18WYSxYy91VF4xXOzSyPXFTKapGzyxqm7Xs9d2Jx9h5YZHW/YsnlXyhLWXR2eFL
WMUaxjrbUYaV/I6mzoPFozTW6DhZPOLSqZvIvdDzo1HEsBf0MhugkGZOsvt4W4FR
2ywAgBatOaLOxzDapwptuwQFeJJL07gM1pGRzCpW/U0M/uo8I5Z7RU76ZATji4QU
QLDVRgG5LnzmHovvfLpQxSIPugWji1ABVy4lJHcQ9YwmLU4J3IFSUnFcJacBRA5y
994ok2givshv0v0+E5hNTiF0iR+HayTMc1OCDpxNYL7EF3L+nMmTLSVkY7veTR/6
7p8CAGbhL6KrbhCUOfwdkYzqj/S65wDSpXkI3yz2swzL0NyJ9KwvnCuDnznzOa33
NZLy2SvWdT0P0Bv8Ogq4OhStHBNdCUVLBjS8r/SSMVd8FkytwgTtgq5/KtNnl3KN
GfRhw8mmzDwU+DDT0FdW6pZykvGwTvyDsMB0412b59ighPeRqI+TQCNkVZLVIxQp
6/BLsWRKNRY3FufuzXCYsGI7BEDA0jOetKryf+blqzVq/jDjJehD1EPfdIEwHhNO
iY/9p+fMjKdoqiLaKu3uKDnAOI3Y64iRFPvihYnrEIkJNXT0hgfyKsHn312ZkR42
5u+xphM2oa/z5INPIc9DCTofhWUvDMQV4QUJv/on2lRBvCU1cvWDL91EKeqoDvei
ZMfgWDXPk9O1RCGCVKszLV3rJgMU1OVKOu2xtiQClD3A0PHEg28xT6aMOYEm0cnc
kWpuoiGxeh5gASskC5oagkseeSYmLXhTlTHzefgjyFoMgysRS7uUymSMzKTYBzVs
itR8nimLwNTVBfJTAYr/3nYWsqyG3F8d/UoF3/W5cV1B9OfBs0CaIG2xVMccL4cO
HFxX9mGPCWQgQ7CKrWijV00gZBlz279evQ18JFjIoPuzBkreE9YFjMaqFxpowOH6
Pr+8yubidnRIG3iz4X1QJ1VW8SS6JMpw7JTVtm6pKvknNh6WEODkNS6PbV8ywy+x
ljvAvyfGiH9wiboOTtIlEHzA8qDOiASgoYPDIv9pwAjhfx/dhGMpNUzFer9NjwIG
+YroWK0k/kw/pbKlxJ8kpxk8MAos6vheWS+5JnWJ8yYPomM8Zb6iSU/pfg8x5NT4
FgCEq4uBCAjXynG+TGRqBZNcZqprUljYgkJluszyCBnuIV5Y9sOaLFaT2N00IUTQ
fa9DunhQBLOZQLKUqRJAcy1gquG/0V6x0Co4NKhck6DZxNU54rYZj9VwcsiFt+PF
KD48Q4JEycqybianrJnMxttnWzoiLYNAFrvjpZmtpsSwKxFHyAiHMnkErNHavZjm
koLWLbfJ5kxMt7LI8XHD2mFtbIWlqj40jJr0wOKXnG3EJnpC0v2mGDdyrDnPAnoM
x3ZUOpSxe8glIDy6DTeVeXsh/wqFFlVq3N1lJ61rvmGfzpZBx2yoGxVHy044qdYg
NbqTjZvArTOwe8SAEc6Go2apXQCRvphvkIL1pHntNs8jJGm5Ycx6CSW5WItjK1Tl
/SiNBMeuCaAPHruypb+FTIvN5kgWax8IbafiMNIwBD7l5ShQVFnX3+qoXzWAVgUZ
NxgaKs64ICnaxuM8jnj8TwIny2WERzxZD60uOaZTF/2rCUj7bKGPP/MknMXe5fBs
HPYPohlFIH9GH4Ybc2KWqYkn/TREnjAbim7G/s2N5b/l+DV0vWFihUNxjISojqcO
gleJC8VKm8wMK6On42BUfCNOgAe9Z+LpUP8mqZLyN+rtjycYVSpfkvmgt7vX2oSZ
TX3YZ5ne4zDJZNlLT0aRl1tVjzC2OL+rqpNGkui0iMXqnKSZVhGgAaUesI3miEQo
GgiMvfn4BL7hhIKRXPUNV8dugaTSrXxFsOKyomdwg6yljVHYnaPr4Eqo7l7B9E0c
EfyotzsRUCx6SddxmbFJcMajgO8V0F4R/SkRH9v9rxVaSsoB+sZyN67KppRcd/AW
gWcxXiHVVabGxdx3mjkpHQ84FTvkSuB/Ggp1sZoEbZoI0XQGyGH5WhHNPCztVxTb
YuVeZDxh5ga67KIaFi3Rtrnn0F51O42a41ZwRVqt/z0V0ENLbGaJOF0y0b/U8IKv
rNuJ3zQStAYZI589Rh9G77RDxY2PoTaVlLVZJqB/cF1XQ+WW8GKKIUpVeko22nVh
M7g26pm6GJXFgw9WxQF2cGpcCHDV6srAQpx5MGvHnfyJF/k7SFjxOajEfwyFJS6t
HsFcjPq2zO81tpLC9tNmmjrLrsZX7qhSgEitAM6zCURtbVI3SIW4rCeogkP9AoWl
EB7Ea5AoVTJ6J5aYQNmTm+DmE+BuPjAqiVj7roz+WYoVrbd5mFR6knu1ltYTP6pT
z1KP/7aYwMgl8jH/GhAR6CGzw/vXmBtkwFhQpkt3hU5X9poNvFV3Gx3+K7st4cMw
J1E6GVcNTeZ2cq4F1d8P3rRIIItYj8pGsC95TVoQ/E4BHRCkyYxDHN0PoNGU1bN1
+vVlQaZHt9LKxy1JSbHz2s3ah8vwcMnzhh6HtWuSSxgYRr/CrPxCjBicNB7C3Gr8
uBf+jJrhwkX0cdj8U7tRTaPLIGtq21kiefLm5V201J/LMaII6vF1L6V7Pumh4M5R
BE12HRO1yNnZfCqQWS3zLbo9C/5FkkrFHrT8/9kRo5NOibLn/BSRi62MU9Enwfma
45vFMkPyxnQ+vk2m4Uh8E2fKmnX58CJa6dX5OXnjl+pTITmwEfKrztCPeDoDl2cj
ZFM4aZdarpdZ7K9VYdb3EPq2mFoJSGSbG5JqddxUyjOLzekuzj4eU2zEajeQ+Ypc
Av3PfgW+je/KFyiwypbja3adkkKLTgmR7Z8DeNoMtXcVrup+lM8KG/SIiZAbJGxE
2hUzAMul4/oHOuxss9bEPioxloxXZvVlZNRvvJVSW6acp0tu7wKrtrxvy0+gfey6
76+9JYas6pZl6Lpgl7TivpdmenYsMtc8rOpl1SAzjyMS0iT09BHIKYyZModaG4PN
+Z7nPPF3ttTHtiaPorlSpEXkyR5wILpV/CuJGPzG0Dggr/TG/bdbwLxk7JJYSwMe
wbU56rD2XahuokPG4LuWuVq6o7n4XO12Kckuae/rMl4CSHbo+6SqYTusV9axAqXW
fB7J8dz5iOSxYkrcE/1rpGYXN/tUKxLFs44cB3oTx5Zv5zatc8E848HeyyS/agWH
Eb9LR/PQYehTAIyJAV/D7BUg0kKYH/FHIDJQDwQWM2wBJLxDl40vlz9zAcsT+h+T
QMpmwGasmtGZwMMCpopE1h0UZ8BtUHgGfHBK+g0EL+LIoMLrQoLtG5Xz3qY0mpNi
RBOEwd8MlVXou5vyYcffhn2WiWjvPMoBLNb2Fh/YIGmQEDTgRx5bmp0GpIyc/nrS
VNf8rlQYBt8PveXGg1+p5EltJoxPIoBfZnR3PeWfCTND/GqcFiFaUJtVc/B5Sb+g
OYN8vhXnawqio+vg03y+io3hBJsXObitTDFzAtPkpNUuCJeKPbDqg1MJfDZsC9aX
qMoGYVue9uAC7r6VqW5Fka89ao1xy3AuK7eonGrZO5iXbBiDjVFGEQZMk5wGu027
WWlTe0V7hWNgbBhTZtik0XUy0PtlPeWS14ngcflTP9ADr++atyBdv45aIfRyNdEP
xycrim/qm0WPJuOaqAaw3erhvxWwUqlpdBURXlh4VNZAMj4qA9l9jFdL1SNgWi7S
w43AkRQsUCVREqTsh9EmTht9fm9Hga82dU99DPwfpxyUotzNAXYB9pyM11ZfLWDw
sYDUvE26jOd0EWtCqOvPc2NowMhuIh0sRruzJijX4aSBLgT5eBkX/Zf9b1GXWGXw
UhyrImTjukgvtics5s/3UPgkjU51ZXdIP5rhvq9okzI9hUpplyoDx7vJ4tELp2or
7RddbTUD3nGuXODeoDjqvLIlKri0cXjcnbyXpvLvyUOkChKdGwKPF17ibd0btjm0
njctw+96Q/aufC+PoMzfJWzXWfuZv8DXd9m7pQbdFQNarwGXu3k4GbMcPxWMjXLN
CIvS5YXbfEIlQ/NtP6SVchu93TgWd3bg/A+3gyiMADPKJ4ccpjdsbhnteETAACUP
yqguL5mC64OH+kGkbDNEQn2lGm/2QZ7Hgp7+EvoTX5pksvAmAbD34uSJeyLYU2cP
t02Ro63fzx7Lchn+t/Q5ZbQb+KP9Mk1Ch+o/zzRdTQ9Bg8u8/YleN4rd8H1rWebv
OpRN+LMFgLumSOZxZX/oAx3+adfzNriOVONtKqnldYzCEC/0z2aeJgvPdMu9VGJq
OTsfmEyF/hUbwn/mUwa1qRBXRcsFUB6Lh07DS4ncUelxTYkkk1dKH5VclxwhBc9J
sgv1m8jyFEo5F4jTgc7m8doCHs2QPyyjQ4cPA3YPW2QjlzSGgWp15HTtG0lPTcuj
g04iDiW/bxnxQUocZFToQA9GnejDZDMBuo58sAvmYMZuVmgw1U1LACkKW5I0b1JS
OBPJXUFYzaKpAKoKppdKnpRq4cv1qnz9jnDmCq9khX8cMVlGGQuhgLT3u7ym2bdU
Zr6UDcBIzq3COmorKO0dMuLVVelEwGKmS1mQFeApAkohgguEthIz+uXK/wYtGU4t
9qaXxGRAgcmQtlZZgn/VqhbCNokXeEoA+/E5TVnmC2AZ9iEh6ozilGUQX7g7Tsvn
yJXmmGoCAZVWfZu0cmDGBTSWSMnx+clUrhOSmyajZhm7Uxo62xtTp2n4QPJ3sPEd
HsdfFDKP7IvLqzHrvdzfKmaZze8gShnvoAqE/XfrZPdWZyLHhBlupNhSotVlcCbt
iplt91oEIwtGFKEi5Asv6esyXcVsrZOpKNhEf3R2Y5LJS2ivbI3jHUWmD8q7UhRQ
CkokwVAnZHCKSJz6JxggBWK5zSnIIrN8XZQPj/X5nsUVK35ncaFBEtOUgTjqO0zF
TtAv5OzZmAF6ZuJNFG/Quq6gOeB5q8mDCD0xYTURLI0GiRCLnGJONoc+6w3sGAF2
gZRWI4+NfQo7wKdlzXENlilohAR5ZcbReKgkQKbqcFmwB0bAJRSP1PpYc7Xc/qQL
jn3TDRCgLYwrWKnL/s9kAXnEX7W3gqaaCNNFZthQI+bljT3O6jszNxiUQ0oSFUvK
hMLPPR/fAH/4ilCo/zMxXsNqzjbdvt3CcK8eO8lIIsHjvVvjPC5yGP0xmLX0cMvG
GDb04aMbo3EFT+/sOmAue9pry4Q8sCagDYbsckwpsgmD3U6lH850Dl3KnZdGF4pv
X7Dke7ClxJbALR8khOOZpSyXXOJQb6w3MMVZaFsDgzj7h0+gG91KKP5QfbCGrrLg
J2Stg7VsbpEFR39JemThA7yWlBCaqsXcZGBi3i4lIA2ONOzF9eSZ7MHA/7XLMrco
dbpBuuhxJ8FP7YqqWa8J0B5n0uFWrVhj2xB0pKi7nmlOvjLTQfP/LoauPoltRafI
iGUwkkrwDPK2AC4q3a/YzDRFcrt6KGc1jBk+WH+t4OAn7k6fkGYsPAirXO3s0WIb
ARKo/r4exibjpUHHAOSqTnXpCo11QWxdtRVt2D4/2QG8rRw2Ydn24oNgOF4nq8H5
kP4n+PhuJrsLcupQEYPPekYLeNSF0sDI8bOxcix8ZX8ORdDboeqaYuQVAVGcULpx
dl7/sjKeVRh3y9thV/F4UfqsmsvGugmuO1ez5BrIyGzf2lGgg1r6b7iIKItC89Lr
ynCzoFFaRUvdk6Ffc0e7cPDBdRRCT3nWEdbuESgNN8DkaldPEuKy6ZMoi7sBSaTM
mqghBeIIV1ANKDLVvcNz5CYCTLP9ohQQH06F5cdHbToy5NvHB1CHlo9dTXS8aYnQ
aQ5MXWQRTqEXbggC2zrra+OXv0PA5u440mEw+7OhD8LxLev6HSUdPaCV1psiSbSG
UB5dnOOGi9a7iV7mwFXI5OiEccVR29ZhHa4r26tSItJ+xC9Kx7DVDN28g4wGkn3F
LzgrpIbdt3AJhz3MDQeW76KsTc/ZmS1stDlMeLPOtnRBOe85hHubGFPvTN4yKgoS
CUVOsTu5cnnIgKoRd+fWrO4OGLWc8dwDloO6lYJieyb585dH8EzDT8HKFvRol84X
b7X9qYwAzVSNMt5AEIxqfEpvTWlICU3Z6solYcu1SFFZnSh75dzMHKbzRn+oE/Bq
uoov4M3mL2fP8eClam9dhSGYf1Icrv+9Dsf36v0TEqlfh0Cm5J6Ai//K09ldmSr0
cB/bpcxYv7PrY3BzLXdWr1J4JXuiE4edb2ETPO1FAdZ4AlWOi4qPhBPFT6H2Yu+e
cND2TeDIFLu9r0kJ4HhW0qANdbNF5GpDENCBVb8zFQM8Oq1uj9uerwdIuh8PHFT5
bqjcV+pivEwZvRK+yFPwiUTWl7Pagy0FVTEscqUvPnd8wUskEbl+RGO8axy3YvsF
qFpJISGMO+BWAXSOPfeVQ5d7Z8Q0YxeD9A673zjEPf/QelwGmDXTmaJC7SA/AQ+g
r0JK51+s/MNLPxplLVTnghGxUPorPi4wB96vcuel0sq19SI5dLkQsQis4Slbb+qw
eLkCxF6bYxFQHfq1FEy7YB9A14fjFZu5ia9YESyB+aULMP2LXquMfTiJfCVkr+6/
2bQY3XijA3kLF/u9UzR7VolV2FK6k1u8wR0ZvrTcAZNnWlVgnZG/5dqp8jvu9TvJ
Vy3kDvSqnsJ+N+kB7LXUPSYtNEhFtJxFyQz5fX/ItG5QBnc2dorHdb3iZsf8hNhx
85qdABr4YneWvEQb56E3tWtGmx3RsXtt0j+7KednOBisizwHwQAiSSuHt9C7C2Bo
GR3LsLnGYcjMO2WvEB0Y+YEcAeQICae+H7Um4VtTgbMd7SZGSnvkdqlMmW9WUJ3J
OY5EqC+9mqNUwDpz9X9Ynt1Im1PW911u76jmu01fk4+KJpXwozQXrVx+lzNBUw5l
sQkY9wBTq4utHs0hRZz5Vj1H2cJuBk+6TBBrA8zSRT6c9rFu7KE4nQmWRMEJHky1
13vKHEvatdo4zTc70xVfzyroqFbHFYb45RpUnrIzzt13pycVP5D8RyigS9LhJozD
YMM01QBf3VKqu1pVfunrgfD0ckAtrk+6jyj4xVFzlUfGyp1g8KB6uVxY3Tx4lo+O
LR/+sAoCHKZAw1kQYBfu8yye7lGkx7bAlSzQlGNzpDG37mzJBRFGSWGiYhLx1YIr
pfPxAqhoTWimfFyDoMBvjLf6SheXWxgiefVWbYaatN7bF4vo8TwBa6x5zmXiC4vy
Llsdu4GYGe8nG25oNtkyOIbvLS2cH20JHQolacOyD9VbQZ69PWTqJrFz/gkeD52t
329tUw18GgtftECq/2CD93YjYwwiDjOp2MGf0xuew3dzjHvsyCiVlvkZjCodUNx+
U/vRk5Ir3TQRBNFSB5Q4vnmpTvd46qmsjPOa4S4l4SLiiagt6SCERJHhoruNdobP
m8l5vkCFdIiA7/8Qxouv/uN9hwSDn0TN6h+P4+mr6nqKWyxIZeBDJCLNV6E7ZH1c
kwM3eFPfvtq0NafuHhnuOP45I58tyzEwn1g8TFpj7696e/K/2HctTZPLnqkgD5fD
PehlI2yNB20T+zLmR0gNzptSDzCleaoc/76hoFtwphHcUgohSrKAa8qYbopyfSEe
mND2SNiJ4fZimQfFUvhNl+tqFpwkfOeQFMN7ETideaFEsQdLfoSSHiYvVlt1Xs2v
+PY9FCg8eWtea2hFa3PuYYOKTEtTtqN9rYiC8HLGtEMpX0IUYr49PRkrPUDE07je
C7uswVRt4cmUpNfqiHrd5dKpeUBR9rK9XUMk+eUi6nB8pTD7W6z4Rh5rW8Hbi8B+
UV0vIzpHOaPwrpRkpmIaCvmKwSJTE/8WVVp/NeMHv/qjncT3hXrg68DTb41BW7SU
ikOwBwhf/OL6pXlTGiVcfqDMy+bKJVefevuSp4qWN9z9gsmFFjDm1qxFIc5yrnOw
A/DDmA6h0kBG4EH69hHmrJ93OALUkTSSVSdggoce/xbf25THfOOb6EzZ0Cr9SPIa
z6dTj5YFQZFZ/zIOV+gBFvknyF30mLpklOXX+e3kdudNGlVG6RBkDbYIDrrrat34
FfXXDSI64dU8zQlecAB9EwjF2Yht0x3+pgCXxv/uzM2O0nL1tb2+XTi1QCV5KIkg
R7UOZHzIDZdOxnlKfSEjCz8uARilapZLv+4xL04H/Y25kjnLEFEe1ATcysZsYEMY
ECko86XOnAaMhg0VHJL5kWG3GWWDbpH2TWfpAk5rBKMJLXecZuhqE0ktGovxdh1X
2Lcs/nk6FtQI0Z6pVHVDQ/n5x2CKIV5WLIvSweIo1om5PZza5vuVQY8Mr6fU1VmM
x3BTgT3v91BJwkCW4DFt8ihWhyYyleNGFqhXriqlPiUsBNSJpoyX+CWyyXyrtxf8
ywHuJWdcAfZvMBrPogFQl8m7NPICmYOzh3zBM5ppRFQiuVSeYODxhUgCIF+Xibyu
C1JoFstqXokh8y/hWwfFun+urIxooNqivIwXwAJSw/34K/+iO/5bJwaFlngDlcfc
WfrTk16QVkgM2YTL2pFhDDtTMrrhz5YG5zJIMmUUxFC49lRXDk9Mp1GNqwsr4yDD
CmBxx0NurwSW7Mga36vLn4uQTj8zfTf4DRvAoj1JCcol30xENRNP0okvijkGf9DS
oacKlkIp/i2bRoE0lJ5tOLC4ZsgpZFXNjy9fNafL9IHXnRjezAHTI9VuAORSjnpd
yhQP5mhHPv79cfGenV/PsxVS6komwePEYlnoctfKLl1s4Koz1dCzDgVKdoNcp4he
bZtdjEFxYJ2R9V3xVAdul0bcofJfMxc3ZNfiFCJcfqijAImT536QRqTaav5+5hqe
bRhZFglphS5wDvRSVI9Bk4CmaNEP0Dq0KOQoPtR0kwPnkq8/iweTj163N/aBK0fH
Ydp+PWmBO/a5CNWM/ZhUYimSg94yPZdPOffutahmFTvsk96ONdsP2n4uVr6Dpo+t
qNQHwl7N4q/2uWwZl3mf8lVIhiWmWFjsxE6/csKKkdTyxPx+QdQ5IlIm4hklccPZ
XgFBovD2F9/fkCHvGcdwCnoQoGDPKsclNa9i2QloXyZuPytwPzhg9qCwsuaWhMCh
iUczxQSV0xr9VuG2ltuNiu/Fg/q401FW80+DGYNHxtmC75wLxDZEtWq0heVvlT0v
7cNgZeJtkDBWl74MrLFP5hge9jm1CsIByUliUvhtbah0BODP8jisgH1NupAeA7V6
qk8PfFJ45gCYfY0rPTapk7Krbm55SEEISlCffoe2z/30fK5fya4AQcHW0xV8uUK7
9VQBSgQT995c0pBcRTYTVGSdFMbbAmUJosv4H1GvEEp0YSiOEFi9PFFS4i5QEW7i
o1gcM9xufSC0XPtL5AKacfZpCn7SqVrS1EUppcMwmkNlZPuqoxbbv+9QgIzgg6sN
Tr6vJDZU09AVBMc5lg+7vcyVVHWLe4hGr5k8t91zKJQqvDuCc+H2p3VJL/9ep+WD
OOWgoVS7356zexCpEKdddywWG+d7qKMYhNGmnc04QZLCAKpTb1SZrRSRUdMTiTWO
hDKsVnxCGXT+EnYkqacgn7ckJO6m8sebQbapK4fZlmcj1yX43M+J6oxFgH2nKFl/
0aGN0Ir4x+r9NnNaXJCfeYrKpeXEab5egOe/4V34IpDlCp9Dkrp0kg9Cfu8dp2Xo
JHt6lhcYBb3uLCIcyeg+9CBpPwV+Db1C/rl7H6F6tSz6LQ2nx3KxThnEFOjvfvRm
5ueSKVLrVF00Pr7N7kyjlcHi5LJNQeqxU/1EnsIdKvAkZZaKmcowGc4xviI+qzk9
gRrXLXRNso0Br75Ha9q4LJtua8ooYg+ZWakypRHFHaXhXPzVnhVv2KhmBMBFzQVG
4nQmfuW/Abr64xIYChGHrp1d5rXdZjv1fAgDYCETQkofdE5K5aCHN2nTmxkASdtU
Ge+uJHOpt6w7Mm4kM38oI+ZaMvIEZ6fFvVgcCPOK4qDqStZz5+f50my8aGYyNCGc
EH1CTfCUhFT95HCKlFgHUNuOY8WfJ3AjQuWk3wpXwHvp+gTXNHBAuOcEGb5kfBMo
hhXPG9BwxZgFTSYp0PQJZe5+MipmP6cU0EOrMqM/enfAI3bTx3A6Cbd90cf4I8/D
at1UVaeOtjO8eFHqtmsIbScrnOr2RgrxKUz77lm4swuPogqHTvNKcJdUvklXWxgg
mxK0YwI2UHtWpdQnH8Do7H845gngIpWTIgBNkdp12vtvTnt4ryR31WWRHfaqw23k
qBNf9MZ8ds33UkIz7ijB6XZqq9z5qrLfqdWWFxprG0/E13hLD8sCIQu/qMtXy0G8
nlI4Q8pLiU/SHab2ugU8+RO53gNmMVW4MP5wP2L589RAuAf5iXp9yEaMgiIZ7Q5c
NzrMtZyWJw45Ham3szcYhe70o1GWwIwXhwZRxrQdXAtTSL7CTZGXq+ffWAATF7CL
ZOJRvazvQclh8ZQ12RhSfa1pX/i5gPQzFz97QgYrl6ZQfn0wz7c5753fixPktG5O
SHm3MRC1W1lfFGlhie5vcD9m1MGnd0M1NO+HG0xUKViR7WuiQHi/pqeDr29L/U4R
Iwm6yJ0LUQPtoTdstRfB0GCJJd3KBQDZ3NaIfSxuSjmaujQu1exsajKd2XBxonlw
GEV01lqOPskcd/pU6t78DeJ85yEKTOG7WSLlul7mY0dKSPjJKON6GqwBhlnR0qgn
9uTc1DdlQZiQ2KCz6tJyt9x6/OGR1P3DPKWdv1h29qEUt3WXPJWJqYQsZjZj4b9E
3SygmfwbzEjxGRyAoP6Cos7rDIQvl8LLT0DywakSfa6VuN+bKYyfkaBIYgRRabI4
PIJfh8TSri3LoiFBFaUKccQU25zc6okY176Cq2XvJDxgdOROLnl8N3rdsKEKvN8v
hxkizIKK7xYwS3bCNocf1y48/TguN0wUQ5IDskfuD/7CTlg3+UoH1sy+60XEducD
o0nqUGiRsZu4fbcRtZsChpzF0cUxEvc0fLhqZ73fzDY6uXTPywTLtmsu9YqTOcAz
mzC00m8TcllliLV0g2/Dbd74Aek+OpSzSjDWMzbCHH+ptq6nnzlWz7T88GQe3kXd
/8iS7LIyuOy5VeCcxTbIkWskjMAP8RMrztdv8kYtusje3RVTIsUi55Okwk2noR6x
lMiTEgR0e56u/soK/X/Vlu37KUov35745DKDEMOLGyZkDnX8YeZLnSPKX/R5L3RK
hPQiLXgWS9Ya+KuCSPmGN4/Ptbgs2KsxpMOE6D5P8frez+CmRUr1xC9rJ3sxNNXB
l6+yIlEPlqsuvza5cy3uz63kFv8JU5+c+ERAPhdCCFtuOMlpx3H42WnaDYxBZhjH
6Zfq5wo2IbxHK5pC9SOglQeZZ7MPK9BNURZLYQxBu708pEr+nTQVFcsgP29LkJPX
A+k9zMGlGI//G/pt2FCNImRU5/3MulZajJ546rABaGrFSTdWapA2krZZCi8KUnSG
xfm3nK542L6b5/spmujktJz9Rza8tf2DjKop27FRcqkmaTFD5juN9sGHNOzkdCzI
GdVeRzyRlyHMfcLnZAclSPP1tuHlZ5qW72/aAk+gXqauhhZI0922WWPkz28AyQ/J
r7OlcxrHHqKT0LQArLn8XHLw1rfpa2Ds+mgD7y7aLOB64MdBYyJ+5MXB/3tlKgbg
6EobGLazJ30vVQVecnnZEq13NvstIZZgXa2ec5QMUy1BDM0xgB5mgCzPxdW6wk7M
QSPIiE6tNypvTaACnYb8jmLLMlPTtsp9RX02LnoPGEBpLbCMczp1cjXaFvvjHGo+
WuzglgLPxjSYexynb+hHg4aglnXEggV8ggq9lLiWTcMksNgSxd5fAH4Bly7UAbeA
ka9voR+ODVahCNgCduzm0Igee0VmKVkFaPkPZVXOZDvsDVBUxCkKMnXaAd8Q9Sgq
oC+13HLr1uaDHFzNz9qjjqMWdlfW5uXUXhaq1esU7LyGtgUyYtZT+v9ifOembfHa
FXEPNbVqPNERQ4XAetBQlezgvwB8NQ9dVifv5JzxBUVv/34nrZb10GfUYVXRT41v
GF/GR+o04s7SwGYHqVtCqrTi/0fz0C3dH2yulSNYX7RJoJNkEk3ZTPaeua3L9zKm
2ngdOcDZ6FIBNblQC+htdLjVA4WV5TMby2qjwK61NF/conHglWb1TkOJES7NLMRT
eQ1oNHd4HREVAhKoWLHau62wiRUcpkL9Xu2/crZUoKtefhlulJpAm3YZZWZG/KnV
pt1cz7kTCX9lG1m+T1lDQKcYrKLQ0qZyV/afch5KvDlnX2haqhCB1hmapSJvE/Xx
sbrMzERk5sWMyIEb1+c4pmF9jPlV/rNTtQBFPBYwCFdo819YFj4XNZGwc/khVDlP
V1eizS3Oscv5peFRjMw4XL+THFO5HMONWq/kiMhL06dqPRiJUSA1giz45ZEYzrC+
ZCtTlb36dh2i/p8IghlUniEGfqp+WquwfbTRHXwdQuDZVzX34/rg2rsSOe2bDALJ
44RY9zfMn6pK1xxlC4ZYTNYNEP3Shk15lYlcdpQc5B6Z6Kbr7IrrI6tWpC+AD+0j
ZmI75hz+lHzi4H03IE3fDe4ecY/evKQ4/DmmbSDM6K2KwwQK0ALdmqsXEEN+UMTk
txlzT0mBwsCgMd/W3Le/LF2VFXSdHqNFs+UO+FdTxWzXUVlZKnpvkBd4d8k3y9/b
+4xYl1kFraD/rTEAqZB1O0QK3bI/OdkMb8ObC8dymAKl5/EGUinsnna4kEtLZqYQ
C2Ape199wAU+FuE3YejEgIGQMFFTPTacsPWFotADv7DzjwWalNHERt4HC1CrdUvX
kcbKAyqDAxvMZURzKerKKsVJzgkMdGHx3EKpK0Ur/SawBYCQNBX/FXk5IY7VKQSh
IsCNFp9vI0F0B9u9nkYcWie/mENkhXE0pusNErh087lKZ+fQBObvui1ZBWpLZDSK
8yEEVz+2e0lvb16JI5ReWIpC2wgQxpQxqc4cYJBYEr2hhOmLJ1Gm5ppHrsuTANCc
3KQ3cywHHAisc1XQysrQ7h2SUFPbq4xeXiOWknQsyiezxIqOzF+Yq0O3CslNj2ex
Z1HBbxD32gb7Snzc2J8+KrbfnXykWAFZwydlwCdEnu838Ft5kk6KqJ2UZXnEyciH
wOFKa8BKPb/gHpGOdeAhu7rJ3C1ggZmpRiGHO/YrBE2RN87JrQPwWd88ddObMZKv
B3elPP9bk2hP21QbjBOABWXLSpYoLwbnwVLKNjpUg40BBGk5yCmRLrVEuewPliHC
8nXcVbzDpr+VppdzFXcHcE50DVKTpokB1x+eWvOiXAitfVsCFbPvDPhA3tq+KG6V
UeeE5yTfrjGneMu/UL9oOoIKpyVzB6S0esAgd5kjPatMWGm74QimBKh4v9WXBLcv
JkekjfGLeF6yIMW3pM8Cfrm+GxtNMPpvMj+YZtmBBQGXwTLdh51tlXrUYsUVNHwk
A2Xap0GFtxtI+jP36d8Z7tE74KGpF44Rb/0QcthQSEwLCsAnano0Im3MOaGs+mnQ
qn0V60In6gB1p522Eue2CvTNmzdm90lB0nYJr2Goc6QFnLj+zQavxVA2gSjiIixT
ISGEZp1dgcxnLacDKCPP8+QxAAnc1BBLVxA3/BMQt7vTrwNLA+kjAUalC6azRydD
82fjIy1qQ48zcepvbhFcxiRg4dBaQiat7mjDOUF3TUI9dtOQqAoKHdkonWgkhrYn
YdEf6OBuEn6PbyUczsjFYxdYc984PoazIL4G6JRWO1x3xW/bywwGgWET14PLIxch
jqaLIQ9g6QXZz2h5q6QQ5y2APDjRzY/HG6zFA/VbJ7+rLnsDge5Vc7s2V0sBIfBg
5vCQAjX8bcZrWo1ZHDzkbYG5MPtFQmNUIKYJZkLsZxK1f59hqdupjijNKJCq0Csl
q05ysi3V+i1WxASmfzI65i+7AGtLN8Y5NcQZttJrcPtRXSH1i6YunW6ZBgjm9l7X
eZGkod6MTP6o5Ffa2COdzDdzapTx0U2T2zuGwWTg0MAUvGqoIpwnxs7B2oGKuvlR
asxicKbjBxcFTa9kPZ+Va4TQfYsKS1qgKBHDajM7Tcqb993h3Qc/B76e21Y0Oltd
bYZrQYxGUOZnTNsQ97j4jHPDAnFAzJiFuXajfdP2APexHeSG3VctPhVuUAowRGzp
2IGGLQm/DHj5UQ/YVpW7dpBx2EYWl3VmVroEI5CeS3LpW2rFHkdbpSzGAjMrpPq7
HH5xaHwlf9cRkZxXn0S8SHP4NeHchPCBEZyB9oV83TjgnR5rMIgHjoX/hMXQOaqx
kjf0MLVgfbigFPkVMevDaVE3Fn0B75M6CuUBOB5lysjEIXTd0VCapf2CT4pnoU/x
kRt/0ICgamm0v1aYPrGwsXQXVIn852bcyBQ1ay27pa3kZS0EWWdfI6+de5Uhrgez
eAdzXDrwM7tWwq8wUUfKrIn6kTufOpJNbuXSYD7C6L2ZbBI2GJLepR5TNIC5T7Cj
XIQVu/xFItUmoQKs7y4s74qE+5xXj6A7aoSlCftWiXlVe3TXm+qb/GrCfJp1zhV4
k/jRIFxVHQrDeZ6D4eWeazDHN6J3ouMXdNCske5LJdU97TwCVPxdAIo5NElrxOyU
IFu7/bVdHIlz4tcjaLvqJIEwyN1xzL+TrJZOk7ejtNcWdFp93P/MCRl3Bj0JdIm2
jnMSo2ff9Xf4GUm6iv2rIm4qkFmI0eGUXBylCja896n00LmjpE7oeae/rWRrhBzm
LaPjR8PRDNQIFERM3d39t3CzJ7KNf6Td14i7iD7T2ZZwhI1HHcvIZas3ONlB9f0i
D/orO9qHBctyu7GeG6RxoUnx+845TaNfV2N+adZ6yvtZlX+0LfsBbxrq9FxJNtUk
WnBfwQhnhdm7qIJnwx7t+DiKpzR6x7skDmokkfVgRV7jZnvnylHDiw448bXZ/qVw
3ma8trPIKkDKtz5eWTBY9DE++ir7l3IG+cuAcFT9XiBRo9Aj5el+NKtY5ATQUrc3
TpDWITwEwWb3ery5XRXzcKZ68g2YBb+kyY35na0FGy40tDqztMuYJen247rji/SR
qzemW7S23H4qYy/S6GkACUQQ3V0Zq2Xclzq0+BmZIL6xew/GVa72LmHYZkko/xQi
oMjPZGe/dUf8qtX2BT6FzkCjgp6DzGSVVI8Rb8Av+kHwKLKKI9tOnShOSegxewtD
hsGKY2xzzZsYCT8z5eWW1mOnl93z+SOHaVhrqqtIY1j7kyrVDrehsJUrg+Ge7LFW
YNRF0r7bomTFvuQ+QlS7hll4Ejp1YEd33mSZzu6VXy8U0vte3M0V0pGtM07wJalb
wdSawcCQn0l1pislU/JEbgdNbB9dPCZpCn5Nrf/KjsWcu3Avg09sB+gPoa6OPXAp
SwygxDdf265bADD0nbVB65GqbuVPKhRcpvGxj5a1TZYpwjQk3UPJ1pUix/Sv1JcA
KfGzjJelvPrPMXdthQAhHKTTGWLvhWgnZ7txsWqZUTchwsldc/cHz1dgRieIV40u
EvpSs0Dkvwz9vgs9zbBs3oH+fR6ZA++Lati8rMgGRt9dWz8UoTBiBHXQtEH2LWiS
qkjqdCxOImXLfcToeS8ahJdkBDSalGGWI4rAIL4DmaBncApTyZ+D3KNZ7hIW73If
0WPpu/kIG8NZS5mofK1URIB5Vn0uzF2pvf6tpOGmQ3Y/ggIzZ/3KqSWNSYnYKdx8
Qb32prKJ59UVbAd0l7YMZWMrUnofJ17HGW7Ts/vC6boamtWg6xOh0rJbyFLUQlu/
NEPIYQwTeOPPpbbD2r+At9EAbVMkz/69tzUVCwoi9qjqi78f4HLCxAl9qerLWc4V
YLOvcLNj4uVC5vbQXLwnPbPWXKgnk1/i+7UiszCCDVljMpNx+g5Q5ygD45ZY6vQU
37Si4BNdxmSwLUZAEZmD+0qTNvOWuGXbdCFOJhjXNfunRk75TI+719uzB5TcLVff
DlTob2jqBlN57x+l8eY34nJ/09Obt+t0KbM5udXeUeXt/cnzOYPDevgrAiDDtX8K
CKreQXhkWMtzUN54vc6s6lOf0jR0+JrbhgGtbtfIFhGF5kJu9zaYKgqonr9KgEGN
d4mDtE2cfVwLbTniVHwZdu0SbbUACRvQEua58znbILQoNmTUy2Ol52xlT7F82WmZ
3nAqtY4yOjFtM4TL2XoVVlyHJ8ZSBZADcBqC0CdUduxu8/uM0eYP2tLxyU7TvAsN
DqHhs6h6iRF+dISl3BHNy/5d8PV7EFWVToDG0hy1lLLigadgNxk9lADP1giiM5RQ
64zoCOLIGBmyAzXB/qOsYkPcdo5w5PSl24uwCpfAzR+CNvu9VI2pla1KMb08JHaa
DSjRUIip2Aq/MkvhB5qM09zmlaS5DhExv6MHzdru6EwOdtZ8H5Fla5x9zxS5waBm
hx9dX2dffkUCBitMdaLRxwzGINz51UzCbc2frL29TEQyuwqHuv4P9gXVi8GJcke2
cYpSjGnVjFEi7QEK++V9MpspAFGv//YKiJ0PADSQSdfmDEXBfalU+KULRDeeYaPt
FHJe7dkj3UdGy4hgGIEYzoEmgeDcasjAwkOwEowP7fD4geGMRVunvJe761Vq/9e6
BOwdujXdqU9Cm/CapfgQyNn5VcACYp7Jpi6LsTEHnDXjQW7BXT7WtFwKFZ7qdutJ
PKCykLZLwIdYOlqqBWGwZvNJH+F1lCaugj06Z1u3oTb5S7rtPRWS4WGoC2HVUQRi
k/XNbMlNSrjnkadn6znb/W4zI7kd2JQqMpxYviHswgUdtMGGjVkWT0kxfZZlg5P8
Fn53yEeDEHoguAsLcqp8LqnBtMeiaK4R58R7AL3MPOl62HqcQWsc3VcbQLVc6lo5
oKIv8FX8YMGGyZTYKMcXNtAdEK94st+S/JpsmIpXG8NOTnL5Q5AFCKtXPwsQYGb3
sdCt1lTGGjkyaB9f2wPkE533244zq83a7+g7wRnMK2tqsHhxXX8T0z+4mU1Ca3Yq
D0rUjtkyVThpD3+OwFEYutmlZXSc5TE4J7tgC5Mf/YJCWr7nmaZ7wtwPBEEf2zCE
vvy6EW7GzFmWQ9Me9KZGsk6n4a+xxQgEEBi/pTSCvPNVIUKmI+muoHlz1eNi1WqJ
R7HxqHJwCClNdoe9Sb7t9Np9VF4+6IYHMlSq+z1l/oob8d8emxGqMj1e5kyCG+TG
w8+YsVkAw2Ill0YNwT7LUXGl4aSgx4CR3CLkEj/VzOsnufEAFDHD6YCy/Z5gMpUW
XjQp8/gCUMcSyZ57kG9r4Jf6SXG4roolZrs2G3THyKqsb96fFzUWbeWjACY3DnQg
unfikne2b6WqY6to0PHOKxMS8frmkOjAXX09E7YtAgoNQR97pRw/hWql99T5E9/9
khKcN23zo7UYQYR/iLQrU5a/KyPkRBMUITc6lSjzcxpXJsUcBT5wa2pEUlfPq5pT
PiO/JHCc/scr3tjYN/T/OIQSf6aWv2p6UEL978LRS/uaG4cJjWU+Q7vowleQuu6o
Q0SVAGJYchybLHP3AE9hMffjM/LrZyl3YexZYniY1w1bTH2NBqQMjhWqG9qmsriM
c6ONeSExCbSQHSPVFusf+3NLCyKPXe3aWQSUY0vcAGVq33dhquI9u6vzSXPeVlxT
1ZH+X031eKw8GOX90aaK2LYL2Q0PVhYmMKAk/5Tc348sbdT9Wv6nh4cfJd9G9czy
NnuZwdjF9OgscHtin5S1HavE1isUSEDhlsl6bNfEXkDs8Qz3tF8YQHrbJs6QT/B/
T+mmUUOE8eQrVvsk7rsWmOTXDULGek4HTJNoMvy4J0BhVjlRBMZ9hG1jLsCkpasE
OE2dDgtHaA7ZLns3fEKtkpeG0f9Ky7ctlzIYP7UmlBN8J8B1cQBZQQWGkXF1er0y
ahcjod4L5evIEy4o0Vctclgbw1imiZ1keAxzUz1pwDsL+qaux3cfzR3PiOVQeiXy
qmTCLJAR6hcaPrQ7v87u+B6iZcLphL1fwc4Kgs6/S7k3yVFqwJCDNe4/VPiBvw8K
5mpkT7JRPrpFa0+WjB2XAvQQJGBraRw2QL69tdoiMHOyPz/ssT/WbW3KEVjg5XqG
2/4OTQaZi7L3RRf5UDB1QBOneW4OY7ZNHcYkNFG0BQokGRc25CFws58FoGfbvfua
kk+hMSgltO1yG+wYhdxTVjn3YnnDwqb/zOtPBoJ0J4Wjjh1A5DWEmLYtdQovZ3R4
5g7q6RnoSmKvPOueQnjsMPxufVhOnvg+vuWLQunqMQLDgiQltLG6lDCRskUBaand
yA+tGFAtzgCWgIX2CpCObxrtlUZtwujkBPoXl8t64ZhLdmMB8MzYOGu/goDXL+wo
/N9j+rdw5pnY7iWZXWESDTEAnm6RCBgi/1WEWxfAsHYSusllfOEWvUiBvxWpGYAr
mthdbtWDXscQO1h5483zxqAbE6Mo0SloWEOIFrOYfdw/lKK3qZnOP3g1aEkJNT2U
51iD3Q+LTWyWWVPF1qjzc+ltxhmnK8edhuRCfAsljOF7CIDs+jOs4d65miJUIVqq
6ld2brdbpLimAyhtwqA/3idp+dRiH2Qps8vdSko7lbxgzl8Qtwnxy9GGMxqOVlQS
r3wxl5OL/4/34cmO6CkmXa+hFeYKWQgBZf8I49raAmf5ZgDDhMsNfoFCaSe4Sv80
ypVj4EC3AtFEEXyUiVMzgulVVlGX4V5EQq0TqVB53wSHo2OMvWTEG8dHm05PwtYN
wjKZCcofLXYqLsUDbjkNTG6Opob58NGxVas868MHxktll7Sp8CILZ/1+r5uZdABH
IgI5SRyWi/0AlBHZARBSdmuAl/zHLzCQYE07lYoz/GvHeNCtnhZEoyouQTJjo2p8
lQnu8UVAdJhWsXYHKMTxOE52jeh/Vivwpi0JJRKpC74i7exrHK9+G6NOrKs7yzNq
s3M/gJm9QkhLaV2DeXsMNFCKeeQjTXqowg2O+tcPsKman/8KfyUr2SM4zhZzd436
HqybmT1DOK/ylOzyz6VVIatUr3Vh6xs1YRze12ZfoBFqHj5TX5LrdPD6p44Jk4rF
+/d/ZL57UAUlD8XgZOV6oIIx+pK9ZJcU4rytEB3mOnEYMV/gNhJDk6VmTRvdc6XN
3ey0mCndmIK19CQlIFL5PClXawtLOm1TNEcHqd4ztiwq0ahb1ArPbkHN1NN46JV3
0oWHCu3zkVRutvXSqbyms0Gas2aQu4AmaLK4BgpTE65G8LFXqJAgrmF9J78bd3l3
Z4c39Pie0Fr4zkYei6mFmEZmpudJPASVNbgDGi0pIKkIVWGBUPM310yWPgiC7HO4
182SgmOB6+IoRasjOSbBoZIiliOOLiZlROrxtpY/ghqg1WBblxu3+tk66kDM8LSY
QxJOh8e8vXUVzGERbXiSg+nA9iYcUruyc7XUujye+iKPOrW6cKVEgoWJHyjGCC/2
SUiifyKI1O0gVuR7eivy5mb/VZqeSI9gUTL1UvfRQla+zax1SrtX9g2N+qFUIRDR
k6W1UEopigU5KrC8TbY7v7wMz3xOQSnWR/l63+4T+anG6/Gm24hXdE4HxGNkakjX
6aIxEcf91XUu8R9btK4JVnbqePTLBU/tyGWFnDw0cfVCz7+AWgqa//JZ6iaEfbmv
alFOuvfT08NAF0FUxdn9z+Rd+dlE8vw1GpNv324ypdvnGOU4WbpRFWCwZesSJUIg
xEZHNWtLgmxNNF8Yby9ylw6rlCQjEZ5irj6bg3OaRYVcJqF2iIU8ZypxoulxO1Ik
+CwaHwEGz7wTRLce4KhFvObNqtocD3rsSm8yBJA8aWbmVz79VNNtNUII43hHU3Aa
+FsLnk2tsq5ZrNLavBcQ0pny/1Lw3iBIs2JmbmVm2Th9NjiB/k0gM2bUd5L8owvT
FMKHZjCrHI+UFmnrFSYWegLkk/ZNBnASisHU9+7Yz5iYg4lx4A5ywnz1G82EDgxp
Ft5jjQtkAIRRaMit0/KEIRp46RuKmzj6BUuZjprKl3+pZej8DEEjm3rEnhW9ZMj0
HZBfpY3A/EIeeJaEdygHXPdxOj6U20HNnWcEsxwTiainbJqRdBVTmiIizHG7Yi/Z
+zlkJPy/r5dX7XJsOkkVddVYKzfeoyLciMgZY10KtJXC2Tq3rcKtF0L7sUVoAHpV
tZFUkq82lcSGi7KdN0/Iupc7EhHeMWVsT1TerpUkEHP+9DIPO5TyBkI2EqOGgUnI
khbpXW0NdMYPfONVpQMDRA9LLaHhvfFhckjSAsyXCkOLPWk/uTJAlW3mD3ef1VzE
vHGTwkY51XV4l7/bomJTtRePes0+mULYahc2zWJbRaup4aqJ2L6Hwqtvp6uYcK5+
r9yA0uPKbKV5S8smPYGzvCWswx6ulRHIonP7l1av8a0AQYlPFD4J6h3tr+lUJuZ9
DIkmPDk0okfV03z0rZg75dJrJ6XTxYBwhdDj4cZ7ytCuGOI4x7D8kOBq6BxTa1Dd
qqGOPdkQE0grV9g6pTW9ZSyNfgXiz7rnrVn4INnIXAkJEd7NHaxkNYfDUUeVUtj6
RVEm+2p2FqxRuyIz/5J1NdIdMO8zgq4Y3Mpxw3DJ64HmyRbqHRjCsL7hURNZ73Xz
ypvN/44sWqOhrSz8I3eeMRj4wesjHaXN1LluN+0AFsJeaW/JgYYPOIjmrkmeZR+2
nfZqxlojPJ8bZ46FEJvWCIcSyBcta2dnOx2yNJpgxQ3hpMmtorQfSUkPjha4sYQ7
Ic6WDE581KXymZ8zPspH0tbT9W55agLH6vt3/eCw0mLNaPf+mzbbjV0W32S0xVrf
uGmTd+gB1lDnvGXVsh89h6dbeANA1UhSUOtgmVXEVTSaCyyvKWZezu2SwLwheh37
gSPbSaVMkR5U2mMVh9qJeFqz32GV1L6fiitGmf9T127fne6QkGt94kpPvQBqkZOz
9nQs98DmQLdn/z+cPD48eW1dkTOJ+WosdEM22JkynaoNbn7jwEguDE4EdeN7UXXK
qY686+6jj5XF4Mp1GZVsQbiGjaHEMtYXSx9mg043uqnBm2DhI5kpGIrIJ6/vXsfs
o+dTvfm4UQmFWtG3KLkukrgxoSqOoAR1CedzOsfqXUN1yq4M3QClmXhh+IhHDnnN
CDvWXBJEXyg45cEfMdetNJORq7Jnl9lvP6qeIOvUuUkYKxe+MjLk8PZSFWgMIRxp
dLBiIYmOYaCUCrxezAhpLplF0UEN1BM/ef7472ya8UarjdMPKIt70BUVc3cyk1XJ
ii2e3HyBEnsu+YUonHO9oQ+8C3VcS+V2zXNYZi8dMKQRjunpf2X74F3ApH0g7Ac6
8kH9BxovldDYXOe5nlj1fvG0SHJFdcyo/IKsGnT5UNfmv5VByoi7LTqCHRq+B0Dz
mZDaeQfcQv/UNeJNPB22JlZgoxBcz15OCQ8QY/D7LpGJoC8qX8Mu/08+fq5NlMOY
wAs71rU7sjti8O49pv+UTi9+zBw6XqswXfhMpOs3kcrfzC7rG1gz8WfkQzoxm+tj
LvRGtYJZ4ZiXjTGazcZKraNuMf2KzpgKpK3XEww2cEPeAqZ73uNkkh4VdAP6FCMx
plWJA4MtPpB5UBa0A/8dJq7acZNBpZg5i1vdIPKP9G1sAYoDgZJh5GREX2Ex3wVy
9Bc7m83sTkpwry62E3/MgldQLmIm0JNfAg3PPmbfN0LIUdOTOTZbWN+nl1lQTaZT
IKvXHmBKwkbFeQmjk+EX8aNZYVbY557qU4DunWQhoHZs743HTea/OOO3ap36bZR2
fMLS1yHQQhqc+C+I55WFrFjeHxxt0D0HP40bwgR1paneTdUpXoE3BeOzz05qwB4L
u4tE94Xs98FuIj/h9Y3626+lqf1y93PNibIce6/W3ZwYOmyli6bjllK2YSQK6+Vy
LlZjsrqAOOpAkPl0kHIuepT39E0QQeEgGoL0jO4vP756mY01nw9kR/XbwwgQqiQf
PpnLLGsfr3c/wtB3846FoTfuO71AyCvjsOFfE+QBeJXVs9o7Gl780aFWBfwy/Uk5
iaDRq+2qdsvwtah+VQk3T+7z3j9xhOgvFC/XZXzcGCxoVF7xdsdoVDZK470vmO6M
RQG9PjsK2dAWYQM5OpDzI5HQ2dfQLFYO7DyBAK5LXAe7SSrs6ppKLE91XJmnjVaA
XKqSyJThkrfMtRtSzt83Kdnf4Y+rVHMHL22AQ138IGh6R+QEBbfLs4E6zqPGvkmB
5yiN0XNiTujwkaqvhac+NWO5stsUqnO0049xjWbhrIrO39AubfO6qJmKthY+Qt0H
N3s7Ek+E+uUI+dem9enFyGxtzCU83U/cOk/BAs3dZbXns1RJqzvmBL/N8T/L3kz+
8D1Vz/L5RCjT2t7MHDrE+UtFmxxj2LB05RTstqOMu1Lx+flJcyvwpuj+/wwO8YRB
Cm8vN6fcgmRc4PHgxyPejKERV3ZHcAfirjL1Q/9JOLlzP/BVry6700E5CoLxplEm
TLNXJEkH2dgaFfl67bMPhsfGZ+amn4q3KpfRUrGSZYccjZOCZjBOAfPg3U6ivJQ7
xyhYVm/wSScQI/zTCgRnPFCYI0K/9ylGr8+//DHsBxf+QX0Qq20dSrUxOrDNUIsl
GRnYa5IWjmPWN3bJ59KeIp7Z7qFEIYS3EnSnilkzdS2KDXvsB/lAlnmOrPTVRX9P
SnpR+2/d39+bYxv3j+VyInj/U8lnutvEF0RFNrPxg+8iXAJGUvYf1XzmbFDidSP6
RW+ldnkgvAPS/y0wcNj1dSXJuQG86P/XLfEcaV9YOEOoPr/IIJmNH3O41NogVsqI
1ST1IvwL2JBgsuHRN+SystjS/rP6o702kSqp5+HeJtoCqRt2/IvbflM5/LhfOxME
AYbXSuSoDDYkoDc2beNdmysGhNFS204KXPCbBW5dNcz88aC3JRWF1JavsQ1ruu+X
a8cIf8os6qNV4HosS8E35iWHAYb9bX+Hfae8ALO9IKSsQpNVSGtbrZ+hFdfs8cyZ
aoV+qhPILfzO0tdlI8FzoNy5B10FUD2/gtxINXmh+IYhrLtDmAH2SWUqrm7N/Fxn
LNtRI4fbLQpapUuVa6RgLkPQzC3rlbo0LKGQD86pNcTPYGLtMKGxyMuA7zNxBueH
x1UF6n+BmAYjBtZJ3i/Cfcft/Ob4vwic/QpKX6NXb1cjoD5Iebev/7ktD5Yq7N17
MfhQSI7OUNtztS44cWgMXe69Ksd/LPj1I90sYVtQx+oc/UM3xEOSEHEwP5IcQBq8
wLpb6uOUWdING+JyE6fzZDAQjKM4XoBtm0ro6aTGe2DbU4E+k46YiImwJCr0+uG5
0W04hm2SBLL2AVAfKhl/ZzSa/vKDRJAc/kuEh6Z1n0mlKDDvZ5uBF8A5T5diwVGz
VWtHf1Cf4DbHM9r+QyUhB2oAlUej4+sXikpLaUkWBV355JhxmIfUERP7pVfiIp0W
IkI8CpVhzCZ1LT0/1sYlpHpnkmvIVmPx/qqwbfyTgGTCbCrRnq0VIEuspklcmynL
OxdYNGqGPQxPaJvu0rNgWJKmnhGA4I2KzsjUm8L7qAwPQZyIOYY6mEVBTV0RPe6D
3CQmnpTcndr6APiQmt50A9ioJsNYDV5QWl7+gl33tzDXIKweENKHcptkLI/flciH
H+t1hy8nXhkmeyBXgNUHfclRYLwUUXE10PZ94MYeZroyD7m0ZK3NPnkWquupg2Qu
aVQZ+blbN1XMGmOPY3vup5ghqsvVqS0M8Ei4m8DVI3oR2kYw9RdNnZpbAy2ax97I
bdLhhuSFCBxb0D8rZT0DOTejNfEdVruZdQcasv4zaOfXYojbo9+v9esLy5E2IVGM
5qCY0PMDvpKKvdGmZymmz19joXuuDt/njVer+vBUbROf5zl12gY5o2ecSK7XEjL1
AATm5azWgyGKdxIsVawoNfNeoHo4YoLYbPjGHUYlD4nt0BWv8ysI6RZII1PTYr1C
Qpbi3llHPsdPD3MEl5oawuzRZ2ISIaSIOtUFvWaBmxbB31CzZ9PArbdZK4tL5fhT
gjCt9nu0FnAMIkCh6MmnS3lyeQv2dLzVHkMhmVQ8TJjgLqBUUhUiKr61Bn0sxFzS
I0Ao+YvI+ohakw7P1ORA0kWbEkrAjRweuxdQ5D9jZlta4464IxW69Y+qRS+bWacb
35XGNiDxiYjEedLRPh88P41itg4QvMAjilLvNYJAEdMnc4zbqcA8aKsSDNLfZbkb
xZaz6ar7pPZOEa1jsEMnBNHJe9OX00aJqng2Hro8H8PjD4NumAYO3IzU290/CH+4
idcx9cC38fFyeTCsdFysGknjcZ6FPNh4uQVbzbvHkk9tD4mdNXk9Wb23Do9FUSgC
Cb9clbrt0dSnDVjinGa0ET0gLTdXuPsvhjTy21oGY2KxfyBOxmcdSRsBNvuwJ94C
Ft8G6KyYVzWZWPIX/DdlaI8GdjDOF5T4xfiToGkusdEA6i4P5kS50meyNjrT+saX
+VkXcvXfa4UIzvCNKDrLgoHWHvpbXo2t4YB00Tp01CdUjjbyzgdDUP1bbQB+outF
Hy3ot2lSCSGDPS+5LrMELtyDkCxPQnsr06iclAteymz8oC4MHsx79cA2sw56u85L
Cijg4HFtWG6/6k7+vOJnuJEG/VoBI5imv2sAaAKpw6Q73A5MPpLPINzbaRYsjfe9
DtuVXm8n0UKAncNHbVfs8ausf1k4Pl1CRuqUsPIGB6u/QCGYU5kjvMBZ9G82iWk5
a5S++i6Mn28BWs33qEI+U3d7GMVaFLeOOWyhlYgKFxXf4yD0xOPtljqKwkGICHPG
/Ns31Eu10e7YC5TOCJ5QYf9Ii8ujV69cwyGOuybF79HctWCwJVMaRHLVOb/zeWTB
//eOijsMBS2O1m5/iXZwCEbJqQb5PoaRM2oBpnZKyFJGCWTU9jo0XBmkMqXllv/L
jB70BbxCp41C8lKTwdmuKdg1rdkNaWnvPw+BRH7xthB25QAlCaEgzL3ja8fHaH17
P2zM0zu/zrnEgxxzhUa/EIzRFcCa3/BrdLjNdm3GCPRKEqW+NFxwlXwp0yJMv5bP
/nb/iWGdosvODfE01Ed/0wVu3i+KsM5ovLxmB3MBTImSdHwqcYG84bAnGJKmleeS
FVB/sEjsxUDtLLpIIBNaZy/TfjI0Oy0f5VIR8eqHYbaUzkGWFpUlud+ictRsgZFX
1UylAy9Ukb4xsMm+kuuqWIX4VIa2IRhidnz78msUvMoQ0JbwXHPqvhGpEt+3SNFf
BuXKyBuADS+oxgu5gruXzZ/mh/OgROSRNEO6BokaUM6a7NiOE/wCC+f/Mjo9iw5G
sM6gCN9vf8OasAixBLPQ/TBR7meBOW470wjWyZXazaxthg/8MlLBrnQVwUnKsz62
vJ8e7IvIKVT6cj+lyKBVgOfYHqMF7oUu2F4T55k2u4rZ3L9mPxenZHEdvGJFPuHt
8ruWCTFKFSoHO+tUSYPZ2UdgL7cPNX91XJOHvQrUh6IXqmN3dW3WZ5EdJt4nLl1/
EPrxQaTqTMeuPX6O6ofmx4BUnRgoKAXckFVLGgY8XZ7SddRruOPHJWzAvW7AV1CH
qjbTO4fwenx624EX9WhIb35I4I8pVybRnrK410ehKyIM1fbwXkych/I+jss06+Ff
dozYg5zoFQF6ps9nDtdbAA7bQzDQ6e/jfPCf3TzDIv18XHrPrBJjx2+9ithhCgKS
65GuuBGljYTKlPPk6Cpo2xHWDBbsk9rON7+mHLZis4O39zPDoUE8kPkFVfbWbMfM
Y6hzHtgaNp8A5xDV/yKtX8yx+2MsWTuGMH03eQrHAwaSWWJIkauVJr28F7WGLKDC
OsLZbKjGhNKCpeNRYIc+TXGET4BlxCma+HNOJjjNLTWCF3GVnyGVo5rXzLQYT6Jo
iI+iTzp078MkQprKywkDqCDFzF/yVztflI8cyQhxq2D//xAWNO9pXV+6N2VvG9TK
eiNTYTXikBO16A5FPsDw84dC1LT/KMbvomgSxY/ngq5vVpIQWD5Do1VbH64HbMgP
xva56+JCcAk86Cn9vh44BNQZtYNsXMxNqMXwVPtAhkOPVGpmiaTh+55OLsXHjF3a
qr4eRk0CC6hnRyQtcGAuzkWRswsR9qBRVUzHN9Pw8NsuyQmX8zDrQ5taGQuRemkS
Co67OwKGpBB7JL5Fb2iUVIbWFAlCFs0ZmGwPMWX0n29vYEHKoHF7wslmibJrj11i
jU9MqhMkMhMQSEzXiDa6fVR1eNs2CTtSj34P2omOlFq2/JI+altl63drNp/WezaQ
9Tv5IJav/7V3cOB244Ay59rrbfQhlyj0X3MrQcumeMtfNVN7DZLOOmrSteUbitnj
SAwx/L4iuiZCPzxyQBegwuB5WBoD6+WnN9pVGbHu8GFpYZv+nd1k/hDSE0aX/14H
/n4cfX7kp4pr5u+46Qhlm16wiCGcCJ9XWjkmELSz85hd+hwE6Oi61wKVDBYIfeeu
J7tOEj9vSplbq9grPVPfIyFws4B6pEb6En2PJdpVm0HVkJ3Mv1p1KImzEBhQFag9
AYKt/CTMZrf0KwxLRDqhaf0H2bzn+dhbg0Hg14+qWMFYfm9wim6gOMiaVPctrUUe
oa6vkLssER8a1rFtL9wac2ZsNSLXjLoik2oXihmPa4eHlc/VhGiV6g7zobShPGOt
z1F1mZNWgvXQbB08Mm21Bg4w42J3rrb2SLRooqlnekw3dTWyitIE8/iMqwyM+45U
qmtsrHLnifdw+VJjS+SoLm6hhoR77nxiZWyI5IviuzfnmkAVZBBdICfRMd8teIs3
EexRWKgBIEDj1j6sPY/NmSscqqVgeylb4X2SSdOdebARtJum8rRSfFDJYZwlA7HO
3rqDry8DWf50LsAUPgtB2sv9ODSefcH4czcEZvoxChXmAhKDL+lmg15y2c5dn6ZR
SPHH90WrF6qv+7mm9W2Rb2BvwVRsh79GApVB0BPno0grqz/24paeWIO3xAEOO2kn
g/HXI1Qah69zLBULc4J+yDiPJOIefoyYbKGVwPgGqttqxKkw+oi/ovTvcYmf5UwD
3nhAvJQl3qsVotEmjEkEzjIvlEGhUA0I/kH8os9D6W1DDaxvTkR01nQVZrfsVqfZ
1v4C7nSc6tJyGw9uHJA1a0J3Gm9tgbq3RIczInNdrJzgb+xhSi6TsTRIvfWMKLsE
eaXZkdGtxRbcdNxQECQjdBU8WNXC+iPCWg0twrpS/MepfAObnNemrEtdOdwIuP8s
+CjVbzz3VPsdLp3C0qu1+rR65K3A2WtnIdk5UAsDV2PV1xBc9MpqGKn3anD5cmNg
0YZrWTJVnKEqMHZW8rDxg1L4esdpUugrcLm2VrXhIVDY3j7eqhaBCU22BHW3KuYb
zTS/5d8JC8j6G/130EoCDS8jsY+a1Fd8bgLDeznIEQUaKfI3PIjoh8NFILHYiIAh
skIIWE/x4keOzduhAuGM5p+9jSqimB98n3GjY9GKVf8TVvVfAzVEGNgH6UzokdeH
U9WEdZ+tW1kWs8JRShLw2lNiemUSd2iSjWXKK4KaBBAjprjHWKqP8KEcGC27BvAd
L4n79z8AsFAKnW8Z+59tkQPyxJdNM0uASbZW5ggb93CxPVN5lA4Q7NpGI1gW15Di
T0+g1t83PZMyuD48h3y+TjUqVhs8O08ou03q9jtC2q6LF0kYQphYycwb2V/Vel3b
AAIuIeCFvTC0PC6vSerkXDi4QFf+5RBbLFAZ+mc+EUL7K3hGx1IKwzN5swRTenod
7+7zxfTeIzKZwcU2oEVcjQYLEGpo/tFbAPLincAKUu6K8vwH+aiGqL6zjHYJv/IJ
fGpzpX/HLi19vCGzh0ptxoBSih3+ks+fbSnBk/9/hMk5IQ/LFWaRJylPzhmFYWUs
DCocnAG1hEwJat7v8nowDFJ4j1tvshcUS/Xa3/iC5Q1XFcMtGvFhY+V322cxdYPL
76kiP5PBYHCnB2gJ42p2MyNh3X1lr1h0o4QT8aTPLHkcQEV4UfUlS3VLcC0Gaq2w
0J6ziFjJYgtbWtTpQJyRm2qc6wcY952qLWJKtbbVhWBBwv+0eVxZLM+c03qI40+1
bC0LXW3Ol6CniGrxIGPMwNBHk1d5gOb3adOgyfCyK32bYUasQLPLZ6KUQv6bEs31
5JNpXtK9Lvb7ZrokALYesymqOQBKnOWzwTtjOA0z6fnk12FGV6221SCdgBXxQytn
NYtTWetVffbseigURJF69NmdwbZL6cHV7omtPR+8L/HYr5VmEpc951yCg5j8MdIR
x5GqimGoCEGGbn1P5zW/TDNmAXo1qxAhLe8ppIJHRICZN0SfEfxEHgxWKqmc5Rt/
xfLqjwN1QmBjJA+lwHkeVdQv8vR2G+JAj/qamfgU3mNeovJD2u9iQCJ7ra30XsER
OHZF2qC6pNISwH9YGMHlH8Mt7O+tQhAGuIbUFvY4lYSO5u/yRhyYE/LsR7BP/huZ
rWHcWnFsbV3ClmY4UslyXc9mmTLcjs5VSvhxEylOK6bEsS/dEuH+LrjftJiINSMm
DGSkdzQPQ/liKsirhYukclrWgUwAUhvwRK+XlYMxtZ6qabqd3LgU7z7jw5KwMck4
D2gIjgMFUg5uUmeN6G77iyCJwuQcPzk3e1TpjPyjjUqacn9DwQj9BPoXGkMOBVm0
p7cxVRXv8qHwYS7c96Ta2yaUL5xqKQw75QgGao+nQP7DADYH0g4gkmKvWbEW6zwJ
4GoFufIpZSduOUpP/VIU6612asYRK91OED6TPNVUkyQ4LDuUe3f9qG9NAB1GD8pk
v5hnfv9Sg8LBLPD2i6Ax77SXhuuPnEfmeo5l6+uwbwdciactFIZOfYUwsQQo3sVP
4xKNql1QSVClRxlI9WTv6BcL/FjTPzQjjDrr/8yxvj4Rj7Q3466TvZEXTi6OF+PX
aVDIsAMW5gJiL1cfj4L/3pIfSEFhpnpDgaZK3UmAFghhNFN4VWbVzKU+9SWj+DQ4
0zWOb9M/O4tv4jGYvPFRuBpfXCfUDXgZ8Ux2oZqSH4m+xxp78mPaNkpI86m/UdSR
3rsi8xuN7I8S7IJDZyEbaaoyz3tVmRivgTCPIQTXHrjxdWdcfa4HPY929H/g4cwA
NQs/hbQF6x+0YnVqqHGkKRoVeEb5hOhPyJKsx2gLWOddcZKclJYc7DbdTnjOBOYS
EkvTpgM8925iTjMC85q9HZ1JDqiQN3vOyrB+Cq7D7g7ye8V//vX5MytngEZi4hOu
NFHVIzQKRF03kdDWZ7ah3dIFi1uAj9kStUPC0OAjv7KfXzCRbY6t6MiDF3DJmhCY
Gpowm0rdXv7ZJlBRPUwVKLVpkwjGe7YAVGirFk2svNEKXF4Us+wkOUQqJ4RNo6yv
2CJJGSOVGXKArmeL4/VSQnE9MfbMNAsZ8ajtrYvGI5j+X4TrwR7q7lu5BM5qInWj
4g/OK7QuJkPsABUkL+p80NBsWCkznyktPE9CIuqm3AddDwMU+DEyXA2kGxpFyHzn
8U4AsDuVcFuTNVpGV2KMUO1F+oQp0LePpMe+7LZTMLWv4xSjMlus2kYjPMfYSAE5
fHwsGHeCSWSEEhOP2z2NEOtk1a/qsUtIUhH/ZgMijy9uDIsKxLqQUY0DPZg8NoDu
LwXCI/Kya3/FVKlhWYBxCQEyYCEtJo4IdAICfPpduqChFN8JpAto7JDulkMsgJZc
ljymRkKZFkuS4QpW2Up7/alfbnL34hW5fXfvG9PeWPfcV5oUMWAPCJU8u/5J+sBg
8XJODp6cTIxLkdpVj+2ushR7MyHWG70PbAIaNd91QpHSsH6kosmULyFalp8ZvguR
uXe8S5JbsYMNCbt8VsiT9H7kxC/k4Cl4QMjm97wGT3zjovFcYNlHEpj2tHCTQBOh
vsdYB2/utPQ8FXV5pghOx2umsXSp88GOR6Y9KPugGYGwgOQIIbYVM4GqL6w/puKt
3Tt/+b+XsGGqOY6HMM7jVKsL+BwrLUg7qt6zbZzrIV+FsZm38AiCBa6E6omyCx0f
C4ekEYKF16TkZ2T57qUFs3aWgQHSR0adnq29qbQAx4jTLiOPnC/aF8sN+lPiAWzA
ICuN2ogvXhj/n7kB4zXc0cEYC8hVg8evDgYz75VNzO76UC1SLaJAzUBmqafOou6I
65ooUZ7sI1UpMdsM5RI89y1Lbdav7hxYhacwkSCRGYekLfbj8oeYdX2JgSFSsRMD
uo/fx5t7nCmozkUqdEXiC1mLzYvvt0ElOveWnVlo74C8vLSRPTqc+wDEKiQpVz8X
owGltuv0GUXCTL7mJR5mXfx+LNL+A0g83ryHVp0QQgasuBE4KMo1tSxVcDuGwtTK
tJAB6GsMi7JHB6I/hIvvMagL9S2EWV+SzZfCfRkfq2I9jzKzN9Q4y52UmkicL/lC
yBn+1iS3eMVAA0oDpO9VHQhEWi8oWbXtrBPowD7Sf7sYfnlGGa/9fkdfhT5M6URf
mn4wfjxeftD/5vyQBvWKiqbgqMoMTvb674C9lPC5Ibr99baXRz5FoMZCOib2Lsim
8vXPghF6EONtH8gg0au1JqfgSBZx5j5ZCDEOk9IOGK/gPUJECkl6NYUQCp69UEaD
mppAR35SchjlY1tUOaZOQ0JyzdR6Ab+QgRapKQS8wu/m/oTD5bCEFNiJm030qhBw
DbHhtMig5qHo2IlTzunxRYu+7Rk2Xk9O3q9a4haxU3XUmzVxZy4S+a0IR54AW+o6
6qn+vJTEO+r3BWdSW6L8xsRg5lUVPWeVVxwS9XzS2v9LCOr0SMwg7MJw7LSkpPXN
0h/8Ml0+WSGzqONuoHH3ZxjL32HGeiDFjb2nxN8CaTbbLmE6R2B5nZQ/+XHLJ6E9
Z0q5r7d8vxUCIGEQSufMuGAbleJkWq1JUAZUNMqUMlphC+AEik8dey9cgqQwPVyG
PIB4P6+o8yeqgzfrKdEjLa05knpn5Z+vOHv6Mviy0GuoUWBEPg/4CUvpIzl6kXLi
7SVclrHtEQmvvmYkcj6qjDhwtYchYctVqf3ks4hfiSmGdbBAFrksToeH7xy4Fj1K
NJITQ+7mvYNhZeFG9MqtNq5inDyMxmaNsxiwrTsn/gPmWnVeDAC+0toFflmdhjhG
Ml2ZALhNQmqwGltux+cLHB8yrSZ65fecirfBte/xBVM7HhNzL1PHhtqwmEYW3fJb
MUca925wW67bla/VBKyLlAXVfmXnt6kstqwaMW34NaoDP68o0HFQWlKByTxBarVt
HEA6rHQxJkh+mZX7mJr5EuPNYnpkv7uhWr0flZLpNL8SDCJ3FBRLwRyib8gt7JVi
/kdzZyHgugILLjf46kKj1S+3xhEIUz/L/SG0/RWDEeEC3ayN3z7vNrfAE+kWfNz7
pqOkZaEWNoFm2wKrkFF+VfXMrgi3RCvnwrsirwKjQYJTb029CH2KhpCko9CiQ+wg
ty6m+UwWiLTyTSyTlfQ2XR28k2tQenlIGh3+QmwTZJq5VryKRKftZ+QAMmOG7H6n
GAOByBlqyJHiDllM7a2m5l1fTofG60pEgX1eeLxXS3RNcRRZ+NUZTxzQTZDXKyxT
Mlhlj7M1rrA3c7eRRY7t9nAfaRnp3TgjkugTkfu7JroXERLjS0yBxgseQdFrlP9v
kDb6qCZ2Uygd46tOZSIhBToKPWxFO2JnplpOs7QlSbZOrq6QMIMjVTZALoy71dxu
iwNMq2yA4xaHjvgvEHyYxBknRdwT5TAZtOdE7l+YkcEpGIUp0deHboqP/12MD4jE
PqNakwLDXmSum4ZZenFSSjBRWPZKUvMGac78acf14i1gWOfzZc/losD8UL19CEHu
ecBZ459XL+/Xz2M0qBM8OcjivVLW3bEFflJxTV6bFY+zBpeXC+Ji/io1GsFUjWDg
6Ov8UXqKtByUUfuYEsi4c4ABJZnHLtH9DfGA8RXq204sRxoZLx5Ki3lD7WRIs2y/
TNFY0TYZpsnI1vqxQpgpIVkx+G/4ZS+95CDDXcVzSpp4U7QkRE4AP7CVAuXoQXSA
QI/4hM7yJSVnyqDzGcG+xSZevbSWs/ojF1hxJDotUCyM9eT2/OLj9uKieKgQPFt8
F/Cpq7ai9/ONOHfDAaZpaUYE6A15h9tLhehugmfm1Ub7etQfF13XuWTt79tTYYyV
89i4kMz/xoQzF7pLxW183Qx9uDPKCEnIPbVqxQLpCb9CwqUfdpvhUoQs3EaHD+lJ
41Fp55UYCPopOMS9J15GmImc7gksiSN6s8mtDfD7MM9wn6P7hSUIzzeniqVFzYRM
OLwYcPH43UNiaShwMbT1Z/HhcwtC9SFHwpUDo+ehZ/yJPyYCMYQu5SYx2aa2uscm
4OYNXTOQkUq1aWBCjtKOjtqRe2S/XEvncqICqQK8cmRM2jzoU2HVudtEZpSMwjsu
U+j6M9OlEU8KZC4nDTfg+kUsH6JIfSj0eJ0bFzhZnGPh2z3dh5v/TmuceC++aL8e
TgFXz2CNn6xOfPZOyB5TSbdwhUxgNEd2AfayferDF+mKS8s4Wrmlkl14ZN9SFiEL
9oCtTyBd+5W+KUNTDsycM1hntaPT5eIhAHIGt8nOIB2/79s+kunSzg3BErFzVNkf
CZyuY0nBwubi/ple2kQxMYrydC2YtUiyoU4O0aEiUeJeApKbkVq2e/vd6BFMNJdR
cMYsiMtLgU5vIHAwKZ0ekHKy6eFIrWtgTQAFm/Plm68BQU/dvy7cAugNR3Z2URvt
cSV+GCEutnS+UwAXbwSlp9NcXL7GQGIDsN7OyJK6MZ5a8t7nD1opbeaTM2xvR3bK
Pu8jVxO0qNLAO/Jix6Ot/uWvX6laTAC4HdonL/ONk39kjAr6uS+n/2kBGnvJIkkA
oBZ3DcN1uadO3hXMkYqxrIl6GDChoyK5LRrmdQj1lzrRl0O7w2gk39UomTerIlDh
G6JHYxSPlncx9OdG5yfw0CJ5bNYCwCQvF2DpjBtv4GCFWr4RXd9Ue/7uoJLD8X4C
CyPgaDVtWtjRQmPBWnbTNHPV5jFszdXF0WcYuAR4icZblyQUxpHcVJRdpXGNsKB3
jRQEbNOlwkhh+Wm9mAgbtWu4WrHj5OTw+lDW4i6Kx7W2OmHs8Z0ElY4i39eGRg9Q
7hG5b2ki3bB9JAzjUZQesXILpLGd+YPxkCqtC+oYs6O0HxuitUjnIuYoLffXcee6
WJRdw2Y3IufZJ7gvj0BxVXbfFv8H0d0qwygwgYlrRH9Kel9RcL8dcfTxAQDdMMTa
74vsgJQAJMJyr1IFDOI0ARQQFdnccfeFKPziQBgMrt+oR8Cb/iwy9PG5MjdkwZ0d
GSvKsQFVVQWvafjaIjlph1spjk/I3SXrjiEaZiPgwseBwbqJMqOJKYvPLsoYMcby
i6C+Q9r4lSusjYtiRPcjPzLVHQZKGXUDeZ/FIpU8mp3VmMxqdvLERkT2Hdcetore
1ksYGYkmmD/fIPxdiLsBbxE8ky9YMuCR9CJGblvkB6xca2Owd199jDQDjSefwF36
pojqFEOSdVrE16alanTlZ013Md6DOEHy/XLR1KniMRZUkPRFZwRyLSaEufFxOn1m
5E5w9pa5sjujAXAUSzP/PyraGaiigMN1l9VLWhILNM958oss38/92WJgAigPDOik
CpDf8bp0okuo2O9nz+lMhQZwp7SCIuzT7jY9CyXatkSQ5IB0hyjSJZRWo1PXR+NN
RxAmT7qRQEBkiWJSlkcsgbeVOGK5nztR3Nexu/p6DEhgvYLxB1XxjsK8efxVNcR7
9xAZ4i+jLRaeLFMf2zIkKAC5oC+OJeEhruhjBqg5Qhwum/NlQ23LIHxAFMB8vU5l
vwAJTOPNXAOUSyj0YRAC5S/WnsxPqr1UU/dsQlDtHIldatHdQKC9Vz5cI2nIz5bz
HMCM8+/yJUDMCYZvEg0QVZCaRVcjyGl7rBFenrZGjVfzcmQ6MaTOXyMg03O5n6xR
JR013OcujbfX4bfFPDRQRPhQ6SshTMp2SVRuYyDCn2BB6M6tiyv0pIkKiTeG18hc
r7IA0Mzk4Ic8YDJGH81mccpBH83oik+co84oPx2ZgA2+zEkOILMEk+3m/Ptkl4fR
7F8wFAbB5rAjKsMN9Wt+UST1kP+lZpj2Ocm33JCVmlTOzyhB9ekmw21rFvfmP4Jj
WrKjDC/faXY4/ScGsVs1Up5kU7gK2Z9AtzYXYlKsf6swmAwO37rtTkxdBc+enZ7Q
1PTdysAOPsQArq5Y6HsU318Y/CvXTAsHdNvv/+2fyq507CrAWBUtnaTDFRWR/HZZ
4RSZPbOu4gKDvsfkEW2hSyb2hBjp7sFGhsUC4d98F6tTgURRUp/Eb/udNtXQHRVv
8ikz+kPUdpzAU9JR8SCWYZlwdDJ1rZlDicmOAYCVfBODcbGVJFeI7cYi/itiyoRd
0fyTjWyLrOQa3DKec5gwXRUo6fhcMgnTTKY1YU9ZTq9P1TUcB0sIlkZ6XJWYdGe7
5gCqOcpXDLUZISE3U4CgI5Y81FlMmesyHFzA2ljp3nhyW0wiy3IB5bZA3UgKeAf0
fRVsTaUtojzXjfw57cerE33iFbkojoGEjY3W5L+yzMO3gyLWGpsv1oLvb5dzkBJ3
ORAEUA2cGzfMbHhU162dDKoltvLPT7InC9bolB2bCR6OwKIW+6vubPFIkFO9LGbR
8aoEfsieHxivs+0VJUJw1GoDuzKJLxx/9sm0QOdqmaaA1NjDmmozvEJe709vGv7b
1KhlhllXglQsnMKLGZgRQWF4s9xxDuQTzT7KPH2cAbnJMq4ig4/JXfQeFIg5GKka
TRJu39IcdaMRFGHMQ3SBfnjs/usBKBAKWnzAFI9pnYMW83byDkeN5gteeE8ujZAQ
dMgBhPavK1++6hfkV+SSfeWyG6Z1ScQdjQ9e7aBLMo/NtwvG84jT78N5FUEvcoz5
SfwAO5iVC3C8PS3IPknG0gDik9tAOKapq11pl1b2PxbpFglA1bQkNTkNLLno6uT2
A0c4gn3n4Tawtoop0+6sJwfNm95fnT60cTvs/Nc/CvY8Y9MXzIlEF8skgEDVQkXf
hWDVMLEw8QWV8BJXjOwbsuzZy4+TDOrch/lR7tv6tP8F/fUEcxB9RCjOTQOaJjGL
WRlrj1Tps+7kOy5ZxysuPNBSDo8SZkSa50MHh1/uC6zAIu2YSHrURppk2m1ceaPu
rPluJx5IWfJ3K+m7YwaxnEUAOnrMJCknBaC1YpjrODBn+nor3/6vTWLp3gHLKFat
UDvp6v3FrKiMXEd5JwDhyULOw69hQvDPEwbMXQQc1Scs9tzA9lcfZlULUj71SOcY
99zhpWP8k6xs0loU4QxzjclsbS27Z3p6xxMCultOzpxaiuEkKPxm47p8HsR6FrDv
BoALOfbPoVC5WhXfhULc8jFS0WdxFItmxok+JeS1JGjDZaJu4eeJTJKQ69sITHzG
kcbzgmOsWwT8cg2FVBtFySURrRuuVbnBtuSGK/L+FKlVbz6PZj4rvy04I3EPFLjW
5AlJ12gpFZaAR+cxDTJqBWB48+cCUi5zc+wadIsHe8AYrjHo+qVS+2ym48QMF9qg
xmB0Y2yiUd8OYQdlBzOm+R2TQV6rxGr7ndBCMx8vkCTQyafQX77c+M2kNb8FVLA0
kGoxXePSkDlGataYFZ2adQeBfeWzDAa58S85z2JV/QfJWIYwjVM9r8H7kSNjQYMz
ffltjrQqczrrUfokuMvBlcfDyyb+yIg+XKUY/QrQia1BC54/TbMcb+hCfSBAgJqn
SBrLdptCcG7QmfkQSNQKdWyrtEqAJJOAMa0QPFTarNyEc65veJtn6UNeoTaUl+1g
gFHhTwbsc2obipUja+RnMjWkwsyBkZ7vrdTk7Xi1vSr2IHHDlvpzmjV4qI9ZqwjJ
/0yVx4EuUlNARitGnAvTBufpOqJ/v1u/1eypOq25jWhEIwLCg+DLaCsbBgtOGxy5
cGiVraoWAj85Ar26oPn9bVTcC2UC36/oyddI+RG2bGwdTajNLGtD/LJ+gpfXniZ6
ui1dHp9MDBJbVcZbyz7+1F60hLT//1lERYfPWe60JI+xvgApV7QsA/p68yPuZz/P
m2Tn2SqyOxT6KZktBTAYU8LLcCUjqNnVbUy3Am/MxyzulAwuFaz2NAR1FvBi8PxT
7uSJscZdYZ3l7mmbVMEIIcsf1YuDvhxDU5RMvMP2sQebWzAFT8AGaensFqiAUc4i
VuJQDBZeQkzfUV1wSbwwEmLNm50XloHCV1dsysO1DKBDK2zRGJn32McIDRldKJUm
p7qfKLdzdUka5/UoM/CEfTRlUcOTaa2o4neKVo2b4pBgQHE4UiZVTFAM83wD5zLx
PxnHb4QqKOmZyW2L5ENYn0BgGQKXPmchDil0ya6Eihi14rikAPDKg9RSPZH6mm6U
OzXa4hMdeD5f7lNOZrPzhViPzrPTJdrhdQvRGMXAmsC0U/aLJr1HS+xIctbIZiLK
Tw3SOfwErdtVQ0Qc/NKljebfs8/K6UMcRZKiV9KmsiOexQ4K5M7OX7ciYgBzb33d
56qo+/iX9L5X8U5F7bTNscTd69wgcMPxVHVLWAYzNdeMC62OqN1uogUP6DGG8RW1
3ZtQEaTCskmqk/sZehL2VxY38LQtYd/WTeDxEjCN5J6RR/AGw22c8V2dg8SFnDKE
xV2S00B3SuGEBHEKLrfle2D0RX/aHn55OGCNQNTKbpzA5t4jkpdjcKhEtwNMP8Cd
pZ42/jNqsPIlufq+nlx1h/IXYuUkCzj3tJ9THcAdSuaSy9WbomWaXW6NhVi8Yj0U
c234rn5i1vqDkk0WGfGRfEkK2d1uGB3tgszIqoLPJo3OlZtZ2FFwwKw5tg2MROf+
H/SzkXhDrKahptJ41GxLkrb+ko001qgqETjtnvu+ex9l+5fyk2xlNzY+xzefUpmT
rEa+AavoMVyHaQ+B5wcAxRjK0ZkY3HRPS0WLUnybETwjLNKRBWCUWxdisdQFt0+M
K7k0gAjIzquf8kKrW9F4eVxrqpDQDJCv4kKpCYkaN0361tvRgTAuCIbFG+s2egW1
nIwWmDIiCo2ci9a6Hwn+Uhw2NlmFx8sv78ZO8BtQk7dCk0gnzp3iUiJoBgkF9f4H
ZWNm/EcjkDF0TUC0AagS9fDscidz2tgaaFAsC50VffU6ym+ziUZTKgyKg+UJGtVB
g2IwJZhix3sYFi9PF658tmIzp/LJ91HqRHSqNuJyg15BI7+GYyUOxsT69BF/oLI4
latF1VM4kZ5G2RI4obY41h6NshcfMdrATFVGAbLGOoTw1tk4usa+6NadyXFtWwkV
ojtHyYDYFwe69cZeckVH9KtyUQ5OjTJT0gaptE5h81s/3FXfgTSCtZRG3F6cKP6i
rnTuBhL1d48kfpxPvqa+Uxy5oKkTo9ggOM/tOjgfWFbphjxlniqtaVBUcpUEC4jr
rAhayf3dIv8nR8vAeYoMnZLbW5d1weDewro4u+0GluZSwhknGmZEtQ6yicmWTRRF
1MfsiCjolLYPTDGTqqlu7SG4OOKXuZ6Gc4bseZ3jb2TefX31FiuvFZHt+9krt0Cp
6xcpD29y8dfhlfmH+2E/rGdz/YOVw5DvM0G9dqyRQ6ohZ9DVtcaRp9st163QYqjB
k5jN9CfAYoCdsyB3Puk96eiFCUn7kdhMvm5u+PJQN11DJ+jKZFN4EfbcHW4XtbEF
IN+J5ccA3kwCWlYHMmk4H9vRkbadV0I9T3aMFA4lg7xDlPxuybIhZAz+qZJy2HSq
cc0QstTxr/gDasflBuEbYKpZMRGMaHLfK9G+h3fEsff8apTi/jExUeahlxX6oXVN
gEexV89n+pg+3lU97Uww95XW6+k2dqytZDHdn/o3MbDLznBqjHCmovbX3KcZYG6M
V199umjnOttOilUivQsZCvIafhinv21rxhuA9RGwMTakU2jxmdjBw6vOn56BkDmW
cALq+GtZ1UPlyYkLh5w2GcF6Pxl7xzgVzKbq+NqKdomeq6+J8jHt7rDrn0BUxSUB
h3vyapmEqdny/hHh53zO2iRzpESlBaXmSf45u2Ws5YBeoJ9iEcnmEZ9BAhyROF/k
QsulpenghoH+rV3w1kBeZolSMAqv5GbpKHDF412nCTg5rdt60OM0WcVhz6AHg9Q2
oXLmcpGcLlaEyAblstlxNMsjcfOz57HFcUtHuHvh9/7tx4KjooXjWr6LTafpBBlv
admn4q7HGn5Q8BnWo3TvxBewioKEeR7Mj94HAlqaIicswbmso6DhujsyG1jCs/Tx
NSeu+bN+G5J1sTNQV63KPKkmHiN05HDw38nVxAWHgA3rrx9zlKIbKu4d2UCVmbUQ
rW+/Ru4dvWk9G3cbN2bDz5hAJBn0LUZxI8QSLdgadigPWLgW8YOpamX75r15Zpxm
/D17/CNi46KrHjdSKjWajuHntSsFt3aPb/pOQtZzRj3CDwhN3vTLktLYAtyhQ/Zx
CQNPAcxTPsGogKRU3iHWej4dZ/I1hvU/44rTMghzTVHcT7asJXkNVFmJkPQTansr
3u0ELIn3UvlmgVKldP0YZ6/akhnFsXAQIC6TH+Ak1rcSEhulmrLKS6Vknx5vdt5N
O3mTdK1Mz1ijN099apZ3anNnjdcwO/gK4WhCXxeVnhKYJVwErHAVe+8nH1ZZ6+CZ
yL46yQ5nkK3QhChbvP0Aq48Ol700DEb/lzO9l6cgWMKUr5U04A3OqrCXdm/iwC59
vknEBVUjHVW3U/hPeKc/qXC80grHQwzeU1TnUcZBFuyn/p6284C7JYbsbkYvjggz
TtQYVycsR1q00QgxAqorFYJOTQTtyr3DvbblQuWKMY7YKT7aYZjH5fIzALU0JKfg
FF4lGiYJ/Bg/DJQi5YFI+X3vW5QZ+mrxGPlttzQwSo40GBZbxvowh6f1n2ry4aYg
K8v/PnmBUkb8v9JSLLeLQjLBPEMSjU1nfOy2WwvMYt3QMqaPm7fiElIjGfkz+vOZ
qecja0MgSb5TcDs9j7Y+TNZ+eFQnCDrvolgpUdqoaBQCMLaZrSedesRma3WkxZLv
/DytgtEqsLuFeEAUh4H4ilwzco9zsiqARPejhaCKzNQk+QSnFvyEhnoIbfsjSJbE
O1A2Lyxy4nbS1CjD+BuCzzzqM1hrNGp3t8Nf79dhaKFcz/V0NGGR+2BzAdg09Evy
n20IawzR6MfrDOSLiJZ26Fqh+AXTSfFGohCtfoBSMFXfo9j8HZqOE6MAjb4fw45+
lOEXY/pN6FQSF1h+lgwt61kopdojOSpa4JFZwBWJx+/IrOB89glAQeNRUOwgL/xF
v+OKSrg7AMbk2d+0i2LK/+0pTcIm9J16q2SmtDRvLlaNOxJ7qUd/dhEwZpGpjrzo
9L5yQKHMqZ4ZWkTE8EL6RUUchOmw6aGzK+eDgiyyjj0E0C7cn/9ziAI0bg6CUAi2
jvx6ltPFktm3QX2MpiWHaB6Dx49mx07Bo5kShshDj9dBlFhfUwIUpFj2PZo0na7p
b/3znS807wlMqbAfwfzEd7V+cWd4RvTPvp8Xp0qpc25mg1bGefx+svh+z8Q1KsI/
ooNu1jAPUYYayl9liSkH+2ocwmxxGY0CE8mhyj5LqMfbXVUdo2xuGcBrIwjbcsjg
s9iqIIXfs1Z8uW4UP6S+Z+/ZFjVf8amr8v0ISNFFXk6MHPZV4THzGlkc/koWlFLC
bWiwWDjPfwyQBF2+2bUvDbuIsyGUuZc0KxOeJ99wD+33AiVUJRzcZ9zzlpKerLYL
RUaezj3RWOn1pu4HlpWVl2k53Ybd4PsKs0XPLPcDQQdr7+oeK3LS9VKxY8aYnG1U
cHWDuYCgcTfXUNe32a5WlW6ZrtlS8zDtGDz+XmNWcJblhnm3bV4yjJ82ozgN6a+C
46Y6ftwh+kkIfewXuXB3zzBDl2/06WmoGz7r1HUEmYOXaOSt3OClOgScbhnRsdI4
UZmsPAr1SXXA4nS4icGXOF2K1quN4uAgXImBm9Dz4j1KKi+4dhXiTGN8k81m6GFp
8ywUEHacsV2IyHAPCuJHGD1c0+dJO9BZydUWGG+LP4gVi7LK1MvhrEN1a3PZegrR
8jdzl1B0ABCO5e32HDADBXhowTehU4lsL2cqjanr7Dwqh0et00pnaSgHW/qnNQRW
lPVaZL7rK+RLKebL8u8sFCQ514sg6On30gseezKTeNlrw6KV03PCyrqt99hr237e
mloRnr0ayX+Iu0cmbKHsO11QFOM8gnodLs1TkQ48xA2S+e+8ZtKNtzxtHYXJk8E+
L3rhUP1aJeZcGrYcu7hcDYLP2RiLm2uV+U+SRv/HeDHqwFtlwg3BSyLN6wRt6bfi
YPcAlQVcQ+6uCp/XPI+RR0bk8U+HchC9DgzmssYK5PSsNR8E6n5xfNsY9BJDOKJL
hDT0zZQnVlqn2T1ODmgKeptg32UW/WcfALWeqR7jnpal/t2a1tbaJ8KZo4IjEqjP
k0093iYxAOh7HpMaudBiCph6GJgdqyGLtXbAwoyWjZnC2lLNlDE4pdlvju6yD45/
TN+wfsCiEW1Cf6fXvrFQpT2gGqBXfNxgn/EhEEkuZkgOvxKDCDqIqQ54axBrGpfD
8Vm5ARsowcpRu0zLs0yY0j5SISjNtEndl5uAnUW1BoFR14fw3P4YemimzX1zR5l9
TvfFISg0rZG45zSIfm2zudwnmpYcX9bTtOW/Ldi/d5rqBaCKaKTqwG1HRhuE3Yq5
BTKkMQH6HkJKz/hOuM88S+oooSawhT3SiacIWGmcc4Lg+lEwvbwiAF6csFxaj6MH
t2uP9HF6AQLG0oA/44uETwB9jiCozGY8NBbvKrRKsZjwpOVMi+7y6ggv0g+bkaCI
ENqYXKRdcuJqrVlpGrkbpJzVo5JMFOy/Q2fBekJuRB7dU4m6QhsAlnOZmExdbNTc
2CUVkhZDU2eP3mVfETvZZkD2N/O+KuavgiLh0idu8gd0EJkqpQBgwPoiKkAuRTOy
PtJkRNRlKkHQnp3UFVoHBq9MMmFkSIBt8LPxbyfI5rAk+CMTw2i+xq0vEbM+0vfS
KLZqH2TNs3Rim7FLzAgKvb1ZpuktL9/mVj4c2EO/fjcwDBYEUc3/+mMSnYSG4a0v
VX6/aVrdiyJHuSUq6IppRGSYcNAa/5UvRJTOTSy3wVodMYBGRlw+W/1v6CLYCcvY
uBpzsA0oK16+dEC/tejncFOPecfYmN+JQ9B6BEUm93iWc1pmfiuREDLuDUbeQVQQ
EAnPS4BSVlLFKtRqb3dZixsrm1LHqBGnjA7oyf9Pj0SjC8N7D5xSiDTDUs8kMc7O
o7Qzvd5+lrMKBFvpDQ9dV7K+pF/+i9I/F8NrSyegZK1H4yUfXdbYk6eK1gYiPB17
XTPu+6QaiTql8xGruZAKwd9+3NBANv9SiUebRfAkreqKlK5iV7nCQZGXI39ExLD4
qyZbhNe7R0gwxxMhxKCUspxYzNTMWxUTT8QxpSaYCS/OYPW9qDC4Ugbg5Xmf8q39
Gp/+thYWt8R4iaxTtsz5hs/Cp02tqFNvtHgQQhXTclF3FBHiahEwC095GeBtpleq
qm2ltKThGvXCECpKgD5WiXskoZeU+BIfNllo3hYkAhtf9g839CUZN6R4e4UX9vqa
9JzJWUhIZJuC/FPz6B9TvScVKdO+Wmzr5BDfTv86YsQfXHHIHHeC+2VvdlGpj2Hn
l2EDQryR+hrNprg0Xm1OsL6HhdGC6h4mbHZCwuEzs85zWGyevJMFKUoIKJnqcxFD
CzQuvAyC4kRjmMrPTY7OJ0+Js//GFdYCr3SuTpj9Y9hkwZYtvRci8Ptj7lJ0cso1
BvjnkivaIgDtJuY1ymLU26gchKkV6pOBWFTJ8OkoDfyFUEMsXAZBqwc2ljswOz2E
56+TDecxbiFNJN8fTnt9eQbWBrnBCMDqwDJ6HprvzWpNCcg8BW1JOyhmuoUjrg7b
4L/6VGlnKdFL+bc+He1SKpb00mYpTrV3yNSkCSSdQUt5VpGYi9YneeIXHtJwCZod
UFQfjgTL/PlFVFpLf4nHL+b8jVfDmFOqFQJ6VNDElqrZJiLIWxUwjmswymcVfm4z
e22CSRFlE2pEKRoKxlCs2RwoWzMSFgrmr3yxFZ80Yx9JaRPm25AFTHR8fbwwORWM
GTj2lRbox77vVX3HCbTq1tGehZuvHYfh+AUgUjVMzVwY+Ub9EoHrnVsLW8EVz3g6
IJ7+dmEzHOQoS45N8fVvMGs6eKbXP26cl5lX/XxiCM9myIdwxzDm5v5xsE00dijm
nOTiMruoa7iF2+UrTub+2YItPkizWRvknfZOJr0+1+wVKa49nk6LICZrX7ZNrumD
u+zxUnU/x6wVgC9CHXcgaT1wofkQCWaxdb6MXIwTw7/zPbYJxmZPmnf4xqjLuQxE
KHutVMEfmIRmzTJ8VzPXexoj60uavjuEp3EgwiAqeJtWN2d4dCeO7saVzfeigJjV
XBpeZ/tlISLJVixzUO3vfDPdtajNpBpyEeCutKifylIRB1ZSKH9K02p4mLQ0kDyq
NReb90+RxHfh/zQrIuszWyVtfHOwns2W+VJ/TiuXBin3ypCEKvVBQQk29cBrDBcc
XBKtAS2V4eyqqFKkahM+9ggNxcrF0dgQv3KaWmkjfwUOZWZD37Rnqci2NxUPdRZx
YbB7QVBHpTRgRzMNCA8tI+uaeK9wnMn1YAZILPPnhrLaGybTILM6sOO4UvVGh5UD
jZ9DgCqB4h6wgBtKPXycxviEHXfTW3CIHvoXL8qpwWMeTM4XQ3Q4cXaJfgOGaMMh
lhmTMPrkPqGIn5ZhVUF5rSWiSd9XVapULJ/VUGxZql7jLtXsI1zAsYjl5F7nCP9q
uLmk0h/6QQKy4SZaEBP6kdqrXo04QH2IKCnuVPlD+2LGvMd+OSHKlzQggv1EafXc
JF4p+EigfszphN0hKIV0RwA8Ld0zai/Mv+KjCiqd77IaJ1xub4NjzNfDXry0ljJ0
Kg080Ti7Y1VjJDYVeXPhRJnu6MmBKxwGAXySGof2b98wUcZsFbRuF6AvfbpRcs/O
lKmaocGpXxiHOuN/wx9zq/ZeFllHRBJsTY4TADoswE3o/VHIxO2Y/AsXlAFM5jeD
qnr/ThZS+icowlFp5x/LAX3jEaT+wjYT4sH37JzKpENwDPVpubLLzfgQG3KoDe41
13MmkpRn1aIA58lc4eOTfEN8deA0oJF92JMB6g2c1xHrMssVzEFuUNMj0bqwFhbT
44DMirb+6AFIFZrqjQpxWuc0FkqLcGpCvisWWzNxXJQ2HtJVC/KA0FFqncz9d1Hx
2OGLezrAQvbG9WdDPLZUr8/kZ8jUzMRHeDpfaWoDzfTjQbpgvTmQJkOAS0hZcyVr
QOu15+RjDXb6qP5UyVTTMc0tumuC7ivsXQp2fCAgOk3riQqIXDjJD+ZBTpkIIITQ
VeWlBD6j7+f2KSBiHzc2wezXYSufaw5VG3xqew0+Xnp0avlr9i85CCxDtOVhLOS0
qW4fW5q93bwCmoHQdAUG2qmNG/wb8MwTbmiB+FafiEYbxGD5nBLF2v+4QoZa0YS2
QFCA8ESwBIAVe0UY0P2EF9yKb5bymGxkhauV52zC/1Ek7iDZPYC6lNU5oaXEhrhf
DqMYQs5rXdsKRBLaWlIf0UyYWwVdKBfVYhkScyIPTI9whTsuGZKhd0HjHdHCXlHH
HI8bcE9wnT9/PG0QzN8oPcsvF3+SpzE3FKeBICQ1vLE0wswWu5zLcwTdfgQ/6VPY
RGxVoYOrkOmH89kGyfan4db+JCiDz4OY1tNZVEs0w0OZlLJ2fh6LyCQofWG/zKGJ
sNqd+1D8y31aZ3emYBXGlaYkrYg2gWddLnCpG8jYDAj9pYEnVFUF7Cnqpff9WF86
6GT/DJo9OJZeJZCGMKt7ktjLvqrqd/dhGv0vl625Qv5+l15wMdQ9iFuDj7sZniBp
pmq4zj98p5ILf1+PfhTbeS89QEukpsx7LioTDWwda6ydH02PWwR7NWiJo4m03OjW
Wd7tSTENtDMcu6CfEgVTrh1T4DYGcCXRAZedSSyIYCSxSbPA6r7SpPhCWyE8sF+P
Kk4wJSmf018Av7amkihNxaalUYkXhy0h2I/M1+su5joowtu/cN0l5VS08fMngcV3
VglwgjTWOdOcw0tjEc3G1flRQT4D7kWebdECN7GxI1ibB7lQKaWYzd5B8sQvIQgn
M0fW5uCu25XqYbdzGVL8uljK+BNpxk/8seVYbmwo2RHObNjpuNwwAL1IkO0NnswL
AvONV31cId7Qg+MI0KXs6JyefT2DFs9y7p+No2mwYwGLZ3+DoBa+WYgxhpdzoYBh
E7xvs28xMBaNfPduc80WIiNoVlNyWcV46V+LO04trhRCL2axvYP/k2FrmkLoHKkD
1pcC1H+to3yx5ao0amDcxC2bhQ2SgpSVVzL9czZLS63Q9j7046/b3G3U0aavcE+M
q/hTrli5/DJhj1dbh6TX2iikwhif9HeFVXQzNW8Vnr+1BbYkgO+XbyHKAdAPKGgJ
5S/N94exofQ3qoV8Z9Cf/U3YQ86Adwywgj3r8CgNtRmjr7PuzXZEyx1TuyUi4wyR
10A/qpu2Yhh9hFX4+gkUi7QcaZgyLF7FxHLQL8/fDtmk0K7gL6G5FW1wyfhtIpMK
ewtKPiOb0IayzaIHOVaW8fGw4vrljE48u+dvvUKweFzaRimksIlkQlTjEt1DPCHE
vrAZfCIOLr+BHH0rzhkNYZ3vIWwgyagP4/1REcmLhsr27XJpvxbGpSnYpSlyxhP8
qis98ID7rTlGoeX35pNRVK2d1Rgi5RfOQ3RLAVMOBN66+bnPoNKy2CYf1c7xHy8H
GFoaGfa8nQNNfxnt4Inx8mkNFmd+baicgOhZEISyAdJQg2jD1EPnTPTw509jzbDQ
pOPRfKt8xPbo+KSOk0PeziBoq/VNOymBsWYoAmK/WcoYRClD9RrRGTjBP8BcsKK9
fM8VrVgFT6Jov/d/id86ZVQ9rXWAcihwo8ii7NAXEqSEtAuqy8ks6EYaQF7C6iqg
inbTwD0nlnQveNhyApL7fsZV4uCgZHZ2F1dfzsYaG1zMICIW9foS6YnxtomcKkWk
+qe/vHrgQSatapIiqiWU96ou78/blx0C5EMXbT0W7q2IN1vmg+wElodSiHBSHI+V
ARdJ464EhRXOz/6jnm+ahEbzhlbmccxC4r6IJmZnRVBictW732sZJROJymTxk8nC
fHZTcyO9IphHpq7yW98Ioxm3NwgMpKXF7XeWfkZuje6ghvQP9BQQbC1TDIqhnmL7
5i2hZ40+5wgklBxp4W2TgQU/ZHUj3Do7fLrdj6Jw5YsGuOZj0xhEpplYOpPpUxNt
M1zDRtGT7GNGjqj+vfQImDp7hcqsUk0I7R5eph3Aj8N+CKS2hhbiJZicTTJ70YK8
AoGUaNkF6dwH9ggB2KkyI/bBbk2rf13KhVC/YDpSmlLCMzMPQvwmsEOOqh9G7JKR
w04JkEtrFwvAgUAuYYNvXfh90fCqVA3d/EfZKf/lLL4F+D6hWhr/oZLOwyzkC4z2
zR+SCejkcNncSfEWRqPJGpp0jJ3izzd5OjC3zycbkd8vBk1CtqmsSsYPawZLkZLD
sCIZDXcmpims4ix5mG3/33ogOT1XhaumYbBEqeUzQiISA2wfBauwmZUdGTc7+RtU
nMKPU197HzUWwsA/DCnztAv4aNkYLb3ioU8tYaId1BNS1PZej1siuoN8jEqqRCnH
+p1IRWMaq+xHON84xErTajkwyjGA/36Fns8v/wizk2EbW9AzV8ivrHbdO903Uz1G
6TtIDqWxDx0TmKvlBGfjmkY8E8S97cbLUumr4iS0n//OqPheJ2G6ZfA/9sie06eR
mBmmFkNQ8lJX54tTLuwA2GRetIJFEFucwQdhcbZzpd344EoKhs6QHBAbXEKS2vSg
K7UKEKMBVhNZdxt3qNhcCzGkfZ1cfbfp3CTzDEFS3CreHoOvt/XLvDYic8h6CPJK
fVLeWZiRInE0SMcxHi8RFZEudacP8rbBdDNvpfSkNKvgmypU34N7aQhg9OouqB28
2Jw2C2UOIwTOpOUAPOHl5LMg34RqwJVUJJU5nfJ+LdPvxi4EnoNEKUlSWhiIMJUr
fpXyyoebF3pFFj8WuFGVB/kH0opoVYTjuM7uMZqKZYAZzXZbDR1fLIRviOFUxvKU
fJysc45s+yPSIjb7fLM4KcKkAY9i43LrqRb7V/3VfuwOUMBBLgvNQgQFRKC3J8uN
nksAKzu38OKG6OJiv5EqcBqdOUKdXn18hl/T+qde2Y6afznUyoUn7H0Gj4wp5dlh
HJb3f3LKLUMQe3AcBgcYYynqKmyz5UStd6rPWQ/TimBKzbB+jyKKdqGUyfm3nFDm
BYabGJ+gRf6VG7Sv7hdm4mi+YILqRhDbUZa/LJrRaliQ94i0x940dC6/P07fng6b
dSFPmAs43HCf2hEkXU62nHI36FPDFm+tpdT84hrDsDAinMS18eZXciHusWWHXJop
F65BL1JI1xdU9PIPgU0kXGN9s6xGRZbV4f+XOGN3S7mJtX8lgR0tZ/dV3nwtX5Dr
3aRtecoQk4APVNeZjEKmG9UhQrwYEzC61T5olz3UOzgHMJTX30tN7OZ5kHD7H3Ee
rFZ1KJwGiRzGmmeQ48OapoXScZALShST4QuJ/bzxR7MxxsSIoRg5RVsEYdOhFn5f
qui7vmhGgsTuNkts0mg1mz/xK2z3wJbm7Zqu498eG/ZMag+Pa9ELiY42x+6kwEwT
ndgcW/OqWaXd8KA9fscitLpyNJfM9wIZ2gH753NcQTznC/1P3iEBr4ztcZqsHW5x
ITc0TyKQeMA1Cwxil42VuJPrMqE311otnJmOm6ub8d9wroniwexd3dlcTj3lHPU3
bk9UCk/UQ9S3dqXMXeaieS758VbzDH8ZEXSKzdGBnP5ygmUhfaNmKzvC1Orzq3qa
A43ZBmTSXbSgFibfX4sEbkmEnbNhTzJnyVAFKZS2QyJD6H384y2rW2nwSzfAVVy/
TPa8aUf6VsUHWYQVfjaRGznJc47IAcRO2047dHet2br2ZL8f4UxFao3boyeUmjA+
DHoyaVgs6xZpxr5qYtgMNv/n30vtVx5HcP5Y9eWGsXR0wHN0FPsW+YgUeCuhMPHL
31HbH0bEnT6soXR90wM3MkcacW05ohNhAu4HpNAWmP7qEJ6MzQ/IJVabIUafp8aL
y4eQjhU1bCVT4XiWMPHgv9esxFNjF4h3x3yj10a2j4F9iVGHLaMGpx92B7tarFec
FoOiYmcS/6sxxSTt5TGUf6W/qdQn++HwRE2NEGdRTWQkt0KpBBqIm5Rukxg2I/nB
+inZV2MOXBVHWS+AMKVTzhkSW87zlaQQM5f5WjDLOGIFLUdmpdNRkHsnetRu5SCi
rxEqzlTKcSiA3wWAxWPC23RTp8Yid20uo9nsA/rfFo6CFOsxk0rwRWTGtTm3XHd0
/83zu0KRsRKOf6Cz5oicV57T+7jqxTPlPgPySLWT08JtXr75cxN2F65XxfaE2OrD
VVLmcTNCt88TLLB227JzHupG3J4VEcwNNnAz1e7XfVu8voRVqxkdjdLU5qIlIrF5
4cO1byK/7RYQ4wQyer1ELN1/eMS9iOlFGXCaF9BpVYzCCjBv27Nip0rAsZktnwD4
JPDGy/fqJgM75uDMw+23woDwr5dk5UASI9tp36txO2XL31V2kEkAKPwjKfFYtMI3
6wIwy4Sf5RFET/DDAPOhBPtg9YpRhDgRkIsvE7eJGXPg1ihRp2QbDMtj3WH2Z206
IIkp8ldzT32YxqRC0vGnKXjh90Ky9jprNzkfMS9vTWYNUem/Nc+PPytPkpvhrUkP
Avzn/6H6UUSZ00/VJ7rrTgy2CoxwvhWU4KiIbYxxeMPPlkr3jCCJOjqA9fU3xYV0
EYyZltTHVIINef701fnPessaxs5mMCkjcdzLx5rpe2NrRksJr0G7gVhsG4uST2Gy
cMq8/EiL6EdT7im8Dgu7SpKBC2J7LjFV8DYotmJc7BYutiSO0MM3F6UGiQfGWhrM
/k4yhqSBLeHqrdL53Tv7cRJkV2XPuQJIof6m9gHeniHQYPsCTUy/ej2ZWjYYhheK
7aLb/3NOLq1agFg3kLKSsgfqgWDD/AoANgJOI4XT4FPumKRxfmkQMp9Wl6R/tDAc
ESgWcdEML136JnJQa+do3izGbvif1tDcHMtxZCPrPVL74KFVdovLkkFeiKAtb+eE
eAhD58mBl+igqQbPxiEGvlCBrpwvNjnL2qoHiKZaf0CxSqCBoAmDKWKyT/ArOlJG
QAlTG9TlWAvU5p7zU96npkc5eADe3AXTg1kf8TkwyHrMLStmVmLBXlFJnpheC9zC
bKbpllHS/c4sZrBlBXzI870jm0ipLdCfojvOOyd01vMxJaArOWzdYhN2EK/C7/bf
rTd2uh1ow3cAmvyUy0bzmCCucMmzlY1sirTckAyij8s9jkb6hD39iuiEDV7zsoEh
r2Og+wtsceGvKG/fJQ8imcZv5cRW6wt1J6XkSfwyKuahhzPhprFcIj8QZuQgUowA
2ucS2LhQSBN6h31tvHuFK9JgsnIMh9oPkfNL3fThP8/oX/OTbk2Qb0y+IwRCwTkR
9guwW9P87YiYIseJIVq0gWxlT5Nwpu8YdQyilqCgyWF+E0vBNC0AXc4bu5e25FUl
HCIgueIyWPI1Cm0XAjpdlZIN07itjL+zeJQ/90gFqX4ViG4ZoIwzFTCkuJmXkLGW
eObVfEqRhz7SJ3Ki55raA9wJaOemDBrS9KRCAQz9QKyMtNhULnm8dSou0AHytKGT
TL/85XIdBjFhTBFBVB6EqEDfpLoBV2uv9mnvATDz10yDBb6Eks30k7Qyyls+vAah
LQ/8SoiNp/JF65/x0Mwx/Rlu3fW750TXK/hpUrdUPvC+jf2HFUqniK1Vu4XXKGZ2
ch+wXwV/JP5WrxULQJa7MFzGPS8+PrcjisQpHpl65Hx8EoLp+IBOPrykK9c2n/2s
Q74EwoVIblGNAp38aqR2dO7ZRxGciHoCTn95WQkjNIULUVrKa2pVHcULaB5GAVfT
e9C8ddomsvS6ysyfD8E260EXqNDkORjucQJwm86Jk+OyQudww/6MFzctE1JT8zda
P85/6ZKtC/uz4PQ4KAa36WE4JXELcn6RFF0Gka2IVXAeyyc8OiBd/63DGLyvdMyf
jcI8wFCq7CF5QxHH7PQQT+6MypAyMTF79/eX16kaDA3CH3LmI3UKmuFTvSeU/COq
J4pVi2jPLy23MJDsqBi9NeezLOqIFEvTWVxW4HlS9H3MOn1fZjD3HgoBD2iSk1E6
JoDJYF92SnXAOYjmsmJrGpYumBUnh1K7/Sf3jay/RR57U8t+iThvYDDElygDBR44
8I4z5jB/LEVAN83vmOCx4TufVO2SAaw5FUYalT0SyPq30V1LfrTdF/foaMc2uPE1
exVic90HYG+ldLVlP/lz6TeFTR23YNZexKFDsE8v/kPmtXfROBP9y1L394WQ5DIl
SVnZao0w8cHgMMA7ecVlAfUwTkZudqEPoLzkOFzqmICbQ7zc9UiKPuN1Ro2FzvYR
uCHXZcuCk3DCh34lAEOpKDHLd7APkM2sfR4PxQ8b3qCwXXK7SrQC8lRh6MWcg3gm
uN+k6jA8zKF1obTHdoLRZ0KVI/RJZ9e/3IHz2T2BSCcFJdgZM/4HLa/WN+wPBgWg
c4wdX6sOO/4+qQViIuqOC4aTRrtsqDvBeaLtDBcWmlX9gmtQHjxg2tgm6jX7lDdS
59QfNSvR7JrqtQy2H15MstxrHhk2+byhqHvremol24ZuWAHueDiR/2u4I3SvZt+t
Wh0RcTl7yKOy7qxc5GCgfcbTwndbm8KcI9S0EHqs1OnMMek9GxRGiIdHW39dY9CW
moU60xgjnvPs+kyo5LWq/oYUGTi1hIUiAjqJQa601W7ENi6xlxxfA+nDBUO/XAYS
XnwL5na1JRTDLSRUviqP5ezSmVyUNBBerPPz5G7+fnf9VA7rawSefgzKS5Jb+kF8
67B7860sxfCuzpBYjaxdr/lCbEVWENEWex0ZPNfrJAhwTpPAOSZShmTdJuqTp6Te
K+CA8Oqp8A8Tz90IEDsgygH5op98cEId0H9exOibJxsV41095upWFtkG43kVIqUb
j+N5ejdgY8IYJfr2uunKjQr7w11sf2kKyHaWj9sn8ubr76/dY57VXp7s7KQvzvbN
Ua0DpesJJtArgWFeXlZ6ySTeDl8JGNBFJ2Wi3mywQPNI9fFRwUS/VZJ0lwl5mBHG
J7XL5qFc4zKZPNn80brqxnCBOnw6MbbdjATGmGkeIz68ifa67QtzgrK3tMIuQN9y
n3LUxJH0tLrH2O1qVc5/asPuL5i3ufW0axzQqoz1+UFBMapN6ekzh9N0g08qVUIC
uXLtffBxGXicAPgaV4I4tMsiXTMeJASMwJ+tYb4cYcy5uaPmrHNDC17Armu2p7zG
+HckdvDCkFRgqtnZxB0NBQ1Ffl8+2ln2J3KESbCrsQdGS4IjLFog8bloigRr+MkA
p3VqfuO0goh/az/9+pldc49wNJNxCANKKezGZuCZSP49t0mfgk+qxfVr+W+5jb5G
hZDoDMh8XrzhryGZ67L+Jq9b1ExYHodZgdUJflswQ182tyorsbbiBuSDKRHMp8Nl
4KxaYThcUheVmKzSSkIeeJyUBb9UDOQ/yElpKl+yn6V5QmaG7zhuMvwsYmrt1QuM
BVczN99Z0RM62EQk1d2Kgn36yLHEoza7sCIkDimkXtmHZtKpVDLxZE6x9NbXLClH
XocYSrNi9lo39opQ68NzRpRgg5NlBFFPAtzAxqN6c41RlZyPfv75+uvCPKLgmtBK
PIummEtLqZUJ6M8f3ii9vZIC7hi0YSNhBqN9inlZpcJBRXgW/hQLCyiyMdHs9wBN
lWLnsO0wf5yFm+1py0f3J57EGljoZunBYGhVFcKoCdSWsGyAzHreb3hoToinw+4g
839GgoYie1pp1tk9DAllUAc2l/b1KX06w4ws0IJi98ZQSU/l/aDDn7ndngXO08ZY
uZilimFk6fXdUv8ADcOxgjkaqb1eivYz2fXs406GMbygFtbb5ImO7BpsYNWzoz4+
pYjGHSO80NyqdhhWMtVlgjVzTw6ENRMUCHt3QvaWeMfDY2amVElJxj+NuehNt91z
jWPKHZQ5wLDOduLDHlhAzioUli3OXS5PyPKgazRaxw4NZtJ8OYiPbwRJeyfVAFza
Hna0Vqv4I/0oMcAdWN2qJmYZ8QQDm7pOzfWG0Rof9qSl9vWqj1GFH0dGj2q9g7DG
dnr97ou1lvbZP/MXZRXyoizsYWZQqE5MWQS1y/c63x3GRujEzFOj4ywxVrdCMSJM
bWbrOKUvAepu8VBe7QtHeMu8E1RnpI8kSVygRdPTGIvyrNFb6NgLZO3UVqXB99RE
dNZTTbAgR6HALcoIVVZjmxvmVMPfYmnWjoXBaQzQkKXh/qsn7JEVvaa0IJhNFd+A
SeLWLoirIb+KwWa9FN5Av5gYFMnRcoLpIFy0XB5wJEqJczxHSb8Wz9+3nIGe+yne
Zm3vgZktDzGhRlpi7Vl7dg9nqFU3t+ZTjD2b61oRstO1JCKB8PJyBCfnAvaJW39E
pwnsyBxAun30iaRNKphKRlnIpXujh0vs6tSlKVk3gBUs55rX86eRhCWlpzeSje2Q
dZ2ODmvApdefzJJeBsvYUUrXcNG7CV4prCdgf5+qxgnStm2odq3hEBuBN7+8comI
+CXKXgg0fZyCcUTsAZLyXUwJ+eiDOl57QthKwFSROVz3H1gxhSzSNXNPK5QtcKi+
/1fRuHQQQel2UP3tJKOIr8dxn8+0dfy2vpNKVgQabPNRNST8Ooz38egZKsxK505V
p0uhEyElojL7M9TN0BHvWBi3zVtKzUel16BVedNJaI+Uept/y/gpmVe+3z08tRrA
PaLM6V8WazAYLhnzrCgbEqAYI8L63Ep9pXdTW6FtLP3BRgNyTfg+bvPDj5OKXaGQ
2mVPpZVzgo0hEeX8QZjVst8NjgeC6n9OwthERxsctMsc0DYE4612BNuXwky9VymH
ETrxLMdAneImFno2wAjaG0fIgHQMLH6tCUlvMmJZ4QJmo3le/iR4HDA/9siw9lAa
3glwbKdh69TiU1oda4OPdcfb965dOK1FcGXg0Ib97R3o3tqtwrDzxQegAvVa3Wlq
+Hl89t7sn4lQaQnBmB1Ediubum7H1175yZoJOUHdo0uIjCRzS/SEOxUzPZOdb8as
/xOEqf7dymbPuYU54ULWJIX0t8wZEnUMNWP4mOi5ghUFGaPah5jd+in5eUgcWg7T
rOqJCen2FukFaAUGDZNXmtaG4M4jPyIPF0dbY0ARx5hfLuXqWMuogH9IPA/DugS2
bXdb66njP4IzitMcP0XttLaPO7NpSOUTpr8aIsP6c3jiuE8udnXB5XXv6h4hSVxI
sv8UL6G3QKY7ob/McVYUsGVZ5zHiZNzm/9Hsf2xk78Z7X3BS+6CEVC73auu/Gz4N
QI7M7rkH20hflb+6ZBxdkvVBYm8JFnV6uigBczxVkCnlI8W+9nYR+RSErSMvs3l3
jwUl/5cutwMGfn9tmrXzOKSieTlQrTMxdJmsFsOcGT7R/IZQ9xOsX3hlvz/guHrv
lcpaOqblNMXSR03oXNXbf7a5rcwyTqaFxoybVdS0cW6WPD3AoIcBfGlF99byzGNb
soTbtKQl2UU9nccY1nduNI/BYbJZOWqJTvcJmu1rrRycsGqR/7NoaEIr9sZeZCFh
hxpXfmJEpy+LS02Tgdp4syX244GYXE9Drog6j6OUGeoHvm/Vk9KfJJZzgNNgoc8Z
7uS1U59/3siLATEuBACdPvStsbRP8iKHaYHerxlYRLzbDOihO6KdwmpuJrTNU5JO
t8IVfQl19rsLre/ilV6JsWOuFAz9D7/swPM2eVuf6g9+jiDviw3jziIb8/A6CW4k
2QnwWsYKL497V+DkhTQySPgtXY90ujzO9cUIsmi2SNo4dBuYv+GR7W/Bz0tVBTap
MNv+gGSeGQMcn8iHoQFtG224SE0MRMjKCDENFL5UjfTMf+FhUn17GxUrDTP7703Z
PTOMvQPu4TcLnm/ZLhILkm+41g6UoJBciuJPbkzpscBUfUCii2v0HBBmH1XaoS16
FatdfXmFI9NiIERUpWIemYyjINNDjo4VjRBa0tNubsNOxdZ1VOtZC7RGT+ZDocUE
2EzeCyFYTwHxec1zfCDtpW0znWNLZBpbULR309meDGGcBk7PC3Z+/8hOsmvYJyt3
OC+PYJl+MmQ3dbNcXGo+0+zDof77EqOlVQY0jj/iKHISsQkmKag9QBC/nUnuEx9e
yDdvVbXeYMki1aOtWRC2ZYePz4cg4UGfnBra+IKtCSn3Q8A+isfwSGyOsZne7kwD
+Z/xw21BeHlXNHNQrPgesy5egWramEkfpvvqcZZakGeY0djJ34jv6zspoKIkRltj
Gjc/E+8aMlZFuWT3Br5P+lyP1L+m31QE94lnhC+FPi9Rpt1Wzm1AxvSc5Cp4Pkex
Y5ggAlhzH1Ofm2BM7mcaAypbI1b2AF67hqv85c6mgkHByX9SR0F2V618MKru8wej
MM0/Qm2CSoNNYoxYrTcMZNmnjiUF1pRVWSb4/HKUUv224HsaAmVd4UfeevUK8gW2
cbb1UHgWDLyVNKJgniWAMch1lldZbG3PGnfKlKgigt+/AstLnOqE7hkaJ5zz/tql
Peyss44DzBT0DEs4LntOCqAY1mGOvzy79KM3KWmzkfl/8BztTuwW+6p577+DEK7x
iF//r6ngcgwUlndGOo8gtdYwlWivRjmTjICLxGqtXFDwxv7YeLLpnfMpxlxG5DPJ
pI0EWyyRNfd9yyRqxrgzMMvjaiiypwrXhW9vJ+yiUPSgYe21nfoRy8SEQNtgwZMB
fXQz5Up/lCOdzcuxGhUohFcZ5UveeE1KHIaWkVSYSSj+KoYyW9nFgJQeciTsWkIs
+mPEmYMmc8skmvyan28ydRaI6bddtYgBDP9b8UIHW1euGauXf54u2i0TwDAvypHt
6z81AYJzFd1xojU/45xKjEAJNfZ1FfLw6Fw/+kPrqOE5DRRfvrFeTUZg7U1bWyCR
4SiKNPMemM0cVG//9wTw0eMsZLGHBPrrBThT0jt7UFoJce/vBUiA7pX2z++J0vFe
d66TU3ns5XOc3o99o09ao3/HAZp6jMp73LnaTcXH7CmQvqGVQui1js/ylKDMbh30
GoLnVdOAiF5asYWuDdJAs5yWCp1inzI6GWd+tOYFhvR208L8ePIHTG2LoNQmSaPT
b+Y0aQvjWAbcLAdGHv8HLK0HGtMms+EpYX14Y4jxNpHfHFTRgCcyN2mLxDhxRRa5
kpGOg5P05qL9mzgTaSXtA/Z0Or/t8Ji48rPz5yjIxwgpJYLcVmQ4Yx9NSjHEB0sf
ZqSYs6NpQEIb4dWiWncW16E4SEwXBDLEL/+AQkW4T3IF6Bz/ymScG9sZSOzkZd2P
7o9Co09+3rShi54lOdHO2Z1twhECAvRxL47KAI7Y4bXrmIOFYPZOLvge9ixbE4CA
cqG+Exgtquo4rg9V+tHlR4pbBQmdldeOf5XAkSw0dN3/LaW4yRPZF5gAWlW2zUJW
wkxIjeb52IylOcDb0g8hPm8nDQJ0wqM86KrNPo0mF634mKVRyfhU6N+yPGDmo6Ze
wZPAJ05R0hN8PutoZBH8v3feGzh4sKdhJzFpKBqw5gmlS0NPpaCFZSn3m4w5kXzX
i32d4bxVaVjozAhq31IbVbq239U7JsutRX5AAIsjQPZ3yET4ADby0maJjDIhdEK0
Ag9gitqZ3k9UQX1S2CJKC9d69Ob/OsXPJdKi/z3cA8nzG69hip9AroWmfSPH25n8
sFytqQtnGims130GL22tf5cYqTeve016bPfaE2KdL9O/khrn5HWCekOjNKoi7DIO
MfXEwTs9gsIbhjRsfouyrjXU2UvKlk2KxJpHo7rFy0v2mD7/ZMz9NN9+FGwQJsOi
3rX9O4mm0hPiD+5dUdn2bcQpAw0E9ySJREYJIl5USPTDZBB53I0u36Z4380OO76W
cQ1wU2bfJvjstYw0gMml1zc0U49SuOPrTjmxOz3ibaX+bWO0kw0YRAKuMWx6ZT+4
cNINmsv0XNp6p3tL+LxnPBkkAMYh5jaKuAVyklykoeIifUgJJzhnqwx5Gv+9GGax
zcc/BCqJRrjp5Xm8SSN6bk/pAxAPRQdYjQE8xQtV4Yy1HAY1QSga+dYV3itb1BFb
AfSC3yTHOanaILIyJz7GGU+vtiPntZEv6Oylm/igOYk2L4s7hNpYrdxruMLXjtN6
r1h0bXGoKGJahfyvCe+Gw6ldbclWoKAGXkIGxRu709f6L4TdrnaO4dF3qclknEkp
e3GhF6CSD61VejOeXBmCRzLrWPOHbS7WYoKtdL6Y7BoIAfBp/qKKpNXWsrN5KJ0y
KxlFnLZzQ4fNZSkudUdtzbaPpsd7mYs8KyDLYBmMtet76GO71qVFPc4M2ITQgyhB
yLpnIlgVaQ0A3912OLs2z+L5FVDuz2RDlVEbomf+G+a/VCAs4YW2vp3OxUaUGWXe
0Rbjf9/HCIVQlYquuTogiJqKMCeQOY7CMkVrbLDj/pWGt3DzXu2mg4s5aV2hZbqI
NyA3LoHDrE6gVqUvdT1FDjc82mkEsADz/pxl4eDG5vNhcatXBx9E4666rR9nuAfy
etj9FZON3Wv0sFGkYiI25JnRkGiA/Wi1rn4oX04O2nxvl43+p3I57q/9Mdxpm1gb
9qzeLlefZglRyBp/rzuHTVgFFVmk/W42P9jNzllfa8HfFcKq20Vo9gVNrCR/FamK
CoKQtp28nU5vhNnIV0UUyg8czLr0Lm6XVQTu5M2jdHgstqEln52HHOrpThXuCvqK
uurhrkWANL4e4RGtXvtXSKfKVTG1HNf2CXYN3/wMDrTs4MZ+zt+mcacaPck0ruXB
pECnkQ4b2G+My0q1KCheZlC3uAevabPumiNrlF66exPEVC63YIz9v9HRxvHE2Rxk
MI3RGuayBxIyYj7RoNG8XdJvYxMX+UJJjCBgmAucTBnlo4XD3yZfd8riRM2Iw9FS
EuA8nS/hgY3c+UWbN/uBx3GZGuxDM2JMfih01Dqn3V1RUwT8T2sbowGMimsKZzjA
Br+t3ARICC6E10z0TliLiiqPk88Ul9XeqO37uzIqXn9vJXRZHR5uHJmMLpmU6KQL
XeN1So6DI0UjnepQNd+6Qwk2sxlt5kQTZkwJZpoWe3cvFjZUJYJs9kAB3Ft6vttr
00RoH1+M4+O2DFrKjUCOUXEQokX1jHrCciR6TNau1/RkCnBpHJygHw/Hjn3oUCRR
QBuhlq0corOGl+czA6VKkWhkdZkHUnlu6ltXHVmw49UVRc1veP6trtAUHksvobMY
2u2MkuLiqw32mEdPjGCfwVFXz1QWyM1iGPdYJsyv/cWqqcsoMrdVVOVTPSKkTPFf
gBGqwVr9gAkQP2b8bo1vowbHl9aZJXJAV61z5G0IqzvVbcFsimXYeRg44msfsv7K
+Qj93AhbfmolyQUAt/GP2Tcr6Svu8M3V06kOvvdDRC0k0AVlmuRaDdWSHZbOA2iy
b8l7WQI404Uo0nyGbVJgR5yng4JaGUl+YSN4YQJfNJ8COd9lr2sv95oAYC/ppzAJ
oBbVH+GMnFVN+wGDx0itQyJ10ASHq7XQ1OsZOJi2gm2hAJqGQDdpezFy7bOqQoP3
Q3c5OYnoSDQZQd2NzWuhmDvR4426uzPhD7TBX1KejoT83wxN7gr/HSzmkFCQZEIe
wt0ZZMEtRTn6KON3VD9pKv7s6M7b45bkoy0SKsYi5HCvcd7cGUViZozBubbJ3cYD
Pgv3iyQ0rfPA/PQ0OVRyj0ar7+RBbG8g6ik8uHznZcaiobTbZSWjx1OxmLunsTub
pfO3Kq74Om5tqVO3r0dDi4OLvHKy8boIbH9qnBRkFdpbwWTPjalRALdXFdOYYOW/
vRsEXz+1sFqHecvYUI8eMOuDdK1ltQN7i/iHZaVRbmTd1xhYlxoGvUwEeAuRNol+
iYYbNLbV8kQPb1BuuOrq4P/kzlHfaxLVZEtqVtCJ48Z0vyncnp9D1UQkxjM4sKGk
GuG8Uc+t1+qGQFqFQoq5svCHwyWqVCy6sOOutF5oy5lmkWtg5q7QA6YwQPKpBXaf
EkBy1czxofIId8pmcrJtb+wN9IFaMmqRDYeBB0SavOW87s8VPUFrY2uuuu6KOekj
ETW43kiGRoU2uLLvssC6U+nokPjxKL+4KOHR0I5RKFH2XPThGBQBFAxSj+mMdGBt
s+sVYuaHBPlUk6k8HLRCiJGFlNCbeLvH/+lN51/IUImchPNCENI4aWtyKVcR5I4c
dczm1dSRE/+mllrW+1WTPPzT5y/iYuJI/umLzw9JUMnTks+0nAlcZkjVzxv0sRZE
QojJfnBPoUoPjWGNXeZ+fbMQkgTD2Dt9inggk+ji9VCpu85+u++knPLtwwl7uhko
0DwY7tL/sSbjdInVih1WJztpeGJPwGbgTos3r9YRXz0ereE4mIaGV6ZTAIgPL6pr
IPNqLLcWtuMuBlrqNRRU2VkTeO+EG0kb6g35RwJ41wnvZb+F9xC9WuUooz684nb8
4iMBitytsEdx3g0wEMz9mvJQPQIVTsHOxaF+oG1ja6obQS9h0hjMaKybiutY8KYG
uTTcJOrVFo45RFgI81BvcDjSieD4LWgISTBqb9Mwhr06LHc7VaZUehkcAHggPFEy
Woz0Otoe22GSGTSTSulDUSb1Ct+1y+MwUOi8m/PN1Tjhj7x6lBL9aLevz38d60Mk
YqJYz9LTRhgeUDGcyzVxnCfIppFnspM2BspCAubGZ+KVtz3Vts7uLLRuxZnzbEJF
cJ+xap9AQjFL1666rMSf9zj484T0R+ULAXdE9Ukzq3ehshi5S3diRXUhWFGkRb3J
1s78/MBaZpYUy5ojqiMopkwiM0OpPlBWNZ842/amwwKh8FXVk8YuICxNv8snDLK9
sAiqnrtRcdrgM+CglIx2D5mj4FdJ3+UqNp2naZArqK3cZ4//RMzaSkqeygd6OxX6
2vSmhW8EUokZb+YA25th5Tn/ycimNey/8UXtsYaE0hbFuwvhltltW6HwIAIkY/4U
fxddhbjBzq7maEjPUe0tJBIPGM9ANlqMgijg7k8iaPN6iFG4ii2zFnWVdp8xwRCk
HTHgGgMH8rk20Jc2Q0DzBC2EsRHPCZS3rW8PTZwo0ooTfn68CRTCJ/dp3lw3dFKO
QnCNzx04+vdhKlX7gJMQU3DjLP+ZbKIlMyPAGWcGABmr1dHVcjuJcbMLkz9pGWZA
OspC62NdyIl/y647nIbgHaf48YmiYzp149aR8ncc4DpnZFnzTKqPzxuXFg1vFbGx
14S9DUxarQs3UbtU5nwBrYvfBVBG1C0oHS0JWNSJOQBA2AX5wpgnfFmO9IPbcsuj
DvIqunuxvZEzjTsmY/1lh6rqfuWQHGsd5ObNiJRGmq6ixFrmIROyL9a6YWrENOpQ
qTy3KEzEzMdMtNCSlGpt4EclOR4mQoD4lt5nzlZrLkG477ReUyFoRwsIdnDoo32C
QmQ454UgilvAzWLwEtQqUlqrCxnJ4bRk9aNKuNK6MCZH4Hwz4OtZAE5SeyUvExLA
9+sEPJph6eDvigCimcNSbKHulZktFMdEupcwRLpuov4aR73ipwoLzudxp48R8a5v
1K47eovv67eXNhx73O22IC5saSuqgBuNWAiZzK565o2kM8MJQYut5vT40XT2wTPD
7BTmmMXiS/o/BQGlVpm6qXfQ+cg6KHZ15aIKQdiod/ExggVpV9ramzbSDThld5Hh
+wcLCUDI0e5KO3PfZMPV4NkVLLbKbUvVWk+PG6atmUcuHVWwv/mE76/rznZyyzut
cwXCMmDxhjfF3LSsWS7otSA/yQ0IMQ3kPbk+Ke4DtxwFUisUGnOOoB6tWLG2TRSm
jVstUNNki8A0JxXHnR4mOhOqVlGp1g+wcRY7syTFLlDeGcXXJKGMmS94Fq9WHtsQ
LhDlZ3d343pK0WzFMZjmb3vZxrw2CcaBhTvg+hlQ78HUx9Mog975IPtl39li4pmk
aryeX5fys2y2AraIxiLLV2wINXt7/2MC/trTMbfT1AbWgEAPx8mj4J9JfGLqxris
xronawOkKt+k+3H+KY31U7w4u7vNjZe72x9kclKnJdS/mop22cQbI8OumRaraNP7
FVUH7lcf9SWjj0jucqSNFtNDJsvHuzoL9RDgGFhzSjy0gnzso9z6tErD6bjumac3
pqg574FgsNDvR3rAUjkp3pmQege5G7fNis+wReGbZ8Xs3XPNmFl9twMrob2hIhNR
zRB+Hwz2dNgCGIPePoHXk0armaNYxMBI+YO9bNrdaUQY1y/n/VzZK4BVOiUbYLt1
sC4nrN6+TB+vR22JJptmjTFhyCJmSjQMrZ6az85RBkS3Zw9d7q4L4Z+Z47W0seBN
Su3TitUs4frlGIiZcWUX+EIkd8A+sIiyAsrJu67JwHPBqX6SkZYbhvr2ZH+WCYrX
yhVJ9FdoQAoEKW2lOG3rLlhzokPE9ND2dJWTxX5Z2G2ihcJMCibL7LuMgb+5aJUm
8bH7WP5HSUgPD56dJjl6ub4IJAHbqim8lua8RNYVfvjoUWptNFW/SDAhsIUn376B
8HkoNjyKWaMtCYf9Hpdsnrka9InAeyWOKTCZn6hyRe+JVRdoROkLpM5AE6LXes+5
Eo1FRvB/85j/kBdXc8vWEEWOdkMRrrP7Lus2z/pm6jQEilV/u4p4CNLHh0KG94oX
dHIQmhf+wG8MO9ywcT+3y2BAijGVKbPwt33ABIi0POFOp+T2FX2lgn1XAnemgwzj
5f+U32MPxuNxftAuu/CSdvUOdHtsDDvCpRLGLQpvAyFCyTKwbV32zFJJ3thWrl83
dOyM84ajJVKsChwR/aUD+ITXWmTyKY1B4o5+/0ceGDTpk5sWNBmGD096bn63x6nU
a+tDUOUZGwYgNuv2JPw0mr8cD3cRBBSDr4MvtvOKcyDNAg8rWcQYJc7zY2RYUUDK
cjX+z+bALH+1+mtzwji6iIIkY4ytwTuCXZdtOGkU1kB/NaxMI+XTJuwmmk9rEgc0
ATD45T5QH4cAz9AJvB7YNmpSCZbJLBo4HFjbKA/A+smW9caTqpmkfnI3WxHJ92WS
/Pbc/yIG3jtoPYMQxB6OgapE6eDigrA2m8Q9j0uuq7Y1fmxhvs53xpwiZ6J4trE7
yJ3+3DuXjIcW6YxklyHMcWvUmt08qeWemrkFTjDf5ngFGebRUHxiyEROxAq8CkPa
r8Of1itzs1TKbAsSk8L0b7JQwcisoBw+EHeqtPtiX2CrjScqo7e2Fstu5yzYIU01
ZA7q7BoofnZJ35NtNd1Qi5wz+70i4R1A4VycImQBlq5Ig3mJ84Vju0Ci0EuLmXXz
uAPszO8qmeUbpaTtAl7A4/0hZkbwHBEmA8iOsTU4D4xXrUBS8W+GZkdrQ/Mh4hWe
4ygqqhMRR2CGGHV7sPCkvf4e8OzoY0M/emTiQfl1uwHwNYWtRjKjzMU+C8Ltwl4x
iZT/Dma1ICFdmfarbCCsBvcgfhTTqWPMheRRj2zDbVrXYdwH/p5pJwuN69uFlyfP
EyitJ9KHetXonxhjzS1iw16XwIiQtYRey8NLSsTo8EJQc6dQEqpHzlpPfC1+xXtA
y3SnwOD7XNyUxGjv0j8Sp2WRE7pBlOJorRubfKBJvPYRagZ2itDkOgM/m01HcaLb
8wqeBmHDdu8O7zWam7QWCsGcNY0hJumTKodnmdlROMOZqSB3wOZq8/fGIz8O6WbP
djhpgC1bv6iyFrrvjl103Td5jax1dcbWVbU3SpwEZa6f+UNKIWRb/wDchwP4hjlw
p6LzQrrM1O21Y79x/TJr3Gz5qfijUm7wxh/fkpjis+XD/mhFeUndPppjvap6zcZJ
0IPm2ysbA+nBERo7D1IO8PnmEbI6jLo0mpeGjobA1gdDGGwzfgBxL1gJjDE5DScC
ILKeSUgksCI9Wvarlsu2Qt/bxNzcrB7M961RJPTFhlNkI2dBjzvSqFBKKYmU6ibz
Jl5ezHtRX6VDxLMIJ5zt8PwXq6X0VylwE6F4vehHiUqPD5hiF1pM9rKO8QolsRct
w7iUU0X9ttl3JeLWKl0tHGUyqNEzSVdTOTeWSGuD/39CtMBsH+T2K2dRqb7wToov
LUBrihIgR7PDkayHOQF6Aej3Ic6y1kDZklyBGfZi03Z+DyAqF/cT2XCiU0S2qYuN
RlvfmhcdZ60ak2ePsgC9G3cgBLiPuWvDQGyOmjGZ8OFb1w0ZLd8Ka8454lUZTx4G
M/7Ag3/JG7Kykv/slEKZGyf1UWcSxhuTSy+DrPU8BYL6tq8G+LD7c4ez+3PIWtYW
TSCzU32qb7xXlL0WqFHfE6swUXyCAmW0Xd+5v4jXQ61TORbEjxhwbM+FtSkuH6y/
TwGqmUxPR7R4kIQi57YHM2l3go4i/Y52A44tlbnBwZ281+OHOsFU0wMWQ5VKCy3v
BGglu3wEOLMqmwpzemKk3qQZF3bZboaJS9qYj8trYr+GZ2/DEB8FlCqmIRoOAxV9
ZNfk16ULYkBpwfzRCKNTdgQuEJfDeRUhvc1fBdBX3soKnr5g/u+CyDeQiboVa2Ej
IFYuan5dPV3UYJU43t4uw8wKnZlOqVuf+/GLViDRJXP/SAx/AgKt66xNmw1Jaos4
fW5dMDzCR5h9N+mK81FeUXaO3IQvCm5OdaOt8518I3YA/dHHh/C6fd3SCFzfUBZt
XnxsD1EAVyRKq7w2CS8ol/uI24qhBiSnXeS8hQCrzmNfK3aUmkaVJB6EyT/klb4l
L2+0P3BvIx/wN4DpQrwUf7qofFif+d+KktMs88egyuQcom73ISMQgIo1KJO3+Nxg
UGko6lcu3XrItHHPaQCGpeZ/KwTWdMsAHq/A8auSp64vU6NzR80OpuO8ncwdxLfw
JhqG5RAqopP0pjksSfD/iI943V7TkXnrWmtF5+wddL6CaP+1aHO4vbxuEigo+opQ
cHDSeXcCXKtP+Bw0feFJZNzfuJnyVHSsOtxIdy/2dnEET7216zsDURdo78uOjRRt
SmseoYq1I6bNmh44Pf03lDakFaFnnRAaXv0edk9cZishroJFgFg7uQ20II6fOjbU
GhJOMjN7vSwkB5LSbrPG5PDmnxS49yKOkUzn8siYAwbHuYHqcf79HdzQlZUnnjAs
SNGz2pQ/38uF+N6JKl4pC0yWD4x9amffWLI4CJ2hEx49M114VsKhzXcirhGHKc88
hEmP+OKXHQpVlpIloygM68q6VcjgryglQlatNbdS3kPz/nHlgmntt/ns/xVdjXq6
Qp8JukYSfbHRNMWpwbs6/ZQGVq0I5KIbGbxfwiiWOVnqGNOadfPSHabbPh2YHn8U
mH8Nhc1H0Yx6CCUY6c42Gf2Hws9s7OnGqgoTedmp9guQuTHWZqoF16x9kniCGBax
ykcs8MhpreYY3U6BDseGj8qC2wS1xhhU8wRu9UOr5GiSjk3EKCaf2q4Zbr1blnPk
+BIvtM+TB6iJaLgHKgksCClLl3r3r4lygE0h1vf40uUfIuLtBDy4zmNzIRBNmQ9Z
T0I9GHEsBHnT0zgg7aRuW2LI7z9SHHPB54KS49tt0rn6VlCQ2jHFQA7Ibt0nnZIV
9TepV8juFoe4yKqGrdpnWn326mksUebizq0A9S++RaBk51liutP9ZUy2oEcbp/sZ
Jx7sKd/bxCtf7pYnpE2u8u/6gEcpf53UAy1FVPWfHmOcrJBn52QVxxgTZDeegk8H
vyzDnFG9rK/T2m9Z2s2ECpzZV3JTlC2jbNQPtXFz8Tgq/yK1zDDGgKfeeaq1QmbV
CE4kSHwLNyANxPp78onafI7j+Ko9IYsAqFxd8casmisxgk+crYQ0iy106nlr+HAh
LzkmeK9hvnsfQ57g4938xe10FGmMqjeIo7hq+jEKpXGjvP1yISqDAW6gtazdvUwZ
OQX4UusA7epOe8ePsHHDvwuwdEW323CjQir454U0KJw3zOtxts1tvgZEnJHSaXOT
8wSop34zw0DAvF8vGpqggaLSrja2u9AUf7AkBnuVD79Zk4l17MlVKV2iu2HPUKy5
5D3uRelJ2ohxpIqID6voPey7XDPyGXlYP6Y6ouf9UAIoxI6bbKDFLwJ5geirMFNs
jdHnq+shCYLWFYH6VjFW7QQmlpZG0UkGjYCDW45oM0bcYk2wdt0PREPe9hMMzGme
ICL1m7Pm4COZEIemUZwZyWkQ5FAOtyJJjHk9Wjy+gFkDLYQ4o+ryK9RfCbg6p4K9
jqpwbfx2JywcZRFRp6c3+dO1whNThtaOs0ixuCWMvj0W8OlLuJpeH4Carlc4teTI
Z67j+YEkscKHbZtYPJWCSYcOWfs1zHdIc1105bdNqOJbbX/6JAC73aZDhEZo+8RU
jnSI8XvqI0/yhBrcHeH2NCrZAFu8h5ZW7d2mVA5i3fjzA+fX69uWFOadJNzagwyV
y/wjNl00O/FNSTDcC2HIRn9nqTMennDv5ZreT386fNNSr4ojlxUdj6YPNO2rl3Ew
bVe7Vt18aZNWQyVyT/RIwRR4yqF7ZyHEmpL61jiGqhgbzgFdz+39p/jhJ5XgQ56B
QHslx9Bxdp6Qp3yCqtbB7T0lZiKh9srC2rlHivmG6wCv8oZhmrmYZFsCXKS0KmF+
AfFXtuCOfMvIjLRG+BPG2ybwHAYz/rnwn38pJ6EEy1/gwCPyitf2R4IBlMGw9xpC
0cxIM5KXEvk6W8eehh0jpMVFFrdmeo2rW7NZ802k7Bye1B8rqIJwRgnezP/D5Nyi
dxscm9J7ZuB9h2vTfY5qJtJDJv10jOTDPwDCyYtCcjNrH/01vvvZKjVXRKiTD9Kh
gUM3LAzo7JkMtgLKc+GEs7bW1g6ikYR/61/7E2ZyaOf8gTixF+C/HnkGgoyqwez+
XNHgOcBW9dZONuigpz5de7CR/VHI/O7AOI1JEhzysIuc52n6yik+Rrcxpo8GlZch
rMqcHXgNlbPbd0MU2Juv6LQul38s+V2ODFTgj9sTO084inh+O4HkcFyt0gdTt629
n4JIieaRjQo/rY3h/4fphaXJfdrXoh4Zl8PiJA0mEren2RVQXExoFUhAMzFBMC4A
8nK85eIgntdUsCkQuIQiGUuDXZ8bMX7ooLOlQMBh//uYwgwx7j+TCErq/zp2ixGH
0cAAyQiSbZWeC74ToOcY0NhWwFFgFMu3whtkdDYxJYcehGgjp2JZGlbc5s+zZAhT
wGqLZg9MZ9HzOWCYhFQljROSe8CURCrs9PKUHzey6LS4/OWtlkjUbMw2VoUFSPEm
39X+KOpwnI0+UhtyYAFpkAEdg0hyCgvWjztQnqs/5dHWw9mFPeOethJviXevNOPf
CD7LmhqJ+GBTyv+5gnkcRfFObCiDZrzMLJa48brHsAa5QkufEajPuS2zB/lPwF7J
pMKQd0m6HK3t0fBqKsFsWYojEVUa0rkdv0VWr9U04AUlK62GFF4jbunx5gcWLKTA
CW3Gi52IUNnsxVjDXMhv59hy9kgK0h9gJiGA2PedAQMQN4aSaZ2byAzspsS2kWV/
i7aSwPD3oweRyxwLW5AalntLy+oQIavxPTXHrMiavbDQ1Ed1Uunb8NdGhe3J4GJb
7ISkWUb8SO0IFnHZMyUxLmLrLJLnBzFwqHTxajUV8uStyDQ12STLuS5pppR4H73O
CeddbptKYT+umSQp2N2vbP0mKWeYMcXhTooWTqPXWC12WOOfAInwv7rLhiJ/llc4
KKPHUF3bqgMfyKkzgVcjckFIE/au9J+XbQPq8TSLwQMSKRcPBKEtQoGib+iiCnQf
JL6tc9uCusG2z+WQNgRgOw4qNiNaLMonKAApFo4kuoqZSSGfsyggJMB5TCGN3m+b
MhKN7jvw9fILOLMRX1wBff2Moo3oQ7ZCNf4REeIqJKGXRKwlFZB8vULsgSDjKp0V
0ZUXANmtQb6qf/KJ2US1lLPbYA8tVWJ7ok3Bo//z/one3Ec29UhN3p20o66+yh7W
eu65rP1boIzNwU/tRnbbxIc0t3JFbPiIDP9GZDKblVgpf2xGoScPW5BNJ/konsDL
/KqS5HWqsFGxHegzSnxLY0tOLGBza0rB5m1QNKcnkqhwlmyiYbLHLrfq3atVSoRK
0diVprIyjCPACfGizgUBjURCamSyBgVb3eBF9iNkWVYNnPRl3v8+SI7bdhEP8/ft
5q7+01HYaVqWAcOgM1/QmTsMdBUlBIXSD6ATBdxfi912p4K3IbbWqimpU1fWCgIq
uTlyW/xoD87NTtwGNaLfE3ApVLSsMzADRnlcWy42ae8hrc4sdDOzb0df8ynHFOF1
vboLMt3N6UGvjKP5jCM/RhII7AoVbqap6XTY0FmLNQwHrE5fdnsuaknnv3yCLFK3
lIwttZr8qzbWDwjj9otAR+Ur2ae46TIJPvchV5xu1PIKRn7z6j8OXhXf4c3rg+j5
tSTMoyV2Ivy7fvLiDzfATOKuViAuZ5DPVpHBAOzsDL1S8OpPn+/J9dXGXUkAdGeA
UM4IcEbASDqnGKICsf0DH771llohJ4YccTBE9omCuxgGZWGA48A+Yyh/nEO96Uy6
G1o9S1MIA2iAbEY3XnLwqgSprMFYgXRGIsCxFe+Q2zNVDPw9U6B/P5//WoYHVE6G
BTkuywlxeN72TQgW9nmqcagQNcVUf+s8jcKRWO/6VHenWPn0BBNeWPM5fCcIfXJl
ikAewMbxpyU0ER+/IErLWAdZAZzjiMHEY+uf/mKQSrYZAwtvgktXovQrjMBYsaVK
RZq3DVEjRxfZoP0LFB74X2YmmYGj3E3W2ayFAlgdYyWbN7BOYe7Us38Zfm+YUEQ8
qENUiVBuRd0ynhQIzvQixKqIoS8B5MTeYYfN12M7BknzxmLxfFU092MQ/HKG2zkf
LCUeMRLV4s8TOWqnHaTHFV7vT3yP6hqvjr8XFuOYIH/Q9F3KoNkQyKITPAJn1Smt
73pYpYO1i9x7AtXCHtx9AUcz47YfUOs/EAWTS4mZVmqow9JBxigEZpwaZI/K8z21
+QcUPK5Ppmf6/+YY3DyNNRaubR1bjdfDzWFp1F6VIDlPdXqaXaE0Y5pCiznTEF2X
v6Lg69v7ZU204ZhEzJVlgO/KjIMMlInb/8MBqP4hBpy1ZbZ7mOwlXrxmr1k53Lba
wnRt4OKlkDepgNyBCrzgRQssmqd5kcfnVNG3rmiy+hvvkzeMBJIkEKdVs4n+HQiA
ZI3g9BCUH2r1vAodX67eSbcGl0MsXB5s1g2bw0ucg/cdMdYC/FGOl8fwCrV609I0
FdLYmTXxqYv9s/igRJGppWZYgVJeN4ZL8xgrngaXcTvJK9CyQeBqdsHZzGeexUPU
cGl3hsuuHlrPMWfdYqMZniV73IMI8c6/WSJlXwtIp8gt9HsMx4SuW3Eeu1CclYS9
HG37/UQqALzngTV5I6WjhSqG33crLD+CmhRd/5JvPr6smWsS4j2IhkZUl9kAFcW6
Ph37WfFaHj+V6A0JmlFVgpAM4uM0r8Vh3apKFiQFzL6SgZ2Ixo+ZLrdR7ZEQL/EX
DKIix1ukE0V0m0j+/sUX39qiWWwteOfI5BbUm/VrA9+QG0MhVj0HSbVooCcCSSaJ
4beY/VN9zJkmjMSFzJNwZ9KBKfCb8XytuhcgT6ix9JjJUE8GkfORtqDG9Ig3wp/t
Z1PK+1QKK0v3Ehz6h7CoQ6YYvPY5v0KVV9jeXpp1p9ukDWHPI2ezMUZ1FcxgQgIN
1p7UHfqtcueieqY7Nj7P0cA1PaKk7ep7H2Gw2NHQAiRanAyAbrLQ/AjC1CcQ7vQd
yVPfUWtxloxZOaDHJu8XvZm5oWRKJvnv5umNdAyC2daOZX2uJ1Gyx7oA20XonAT3
fs59nD9Q44XGqA52MBRw5rBHDJoVHAdSPLH4pkI6A1BQSk3+ywWYJov46AS8PrAR
NwxsePsjBjqDvx91J4gLiJPnbbaJZPRvh6mKu1lMYebt7MmMeMViF06suO4apKad
fSVdiAMW0FXIIa8VFtZQSBPfKlIa9NWEoSVRJ0femsK9qt9IokaKe87JOPsI7wDc
xfG6UBExMxz0F/yld03BEBXtbkhGn7hJIUO6LJisws0vjV/XCU3BhkmqyNBz0Cd7
hcebe+XnYDdwiRtEv767OKlwvj4pBIOF9EAfherDaHYYeP5e8yxABiWjrcHt987e
OWXyzULIwYU/5XDP69m6Z/diyTgVtbO24MYJyVpaEfD+VYMYinAc843m0s5owC9S
BOdWptuZja94lJzRPXAcH97sZi3d0rVNNpExjr4K4IhpWHx0Pah4JAu89iufYP5Z
FGpGKvTuBPSAaf89aE8jE3EJbxD4b8wtDYAdf0SKf6q5SZhaDTrD3I2SswCMwt42
qClF7kzgktpOeCtVWFKL0ruEKOTlxL/UT7zksavdqGpl0SW0AYdhlRJc+pT535tS
qsKLxCU6uGv3efihMsYSJoTezDMlcnJbHgq4xXm97Nj+NqHHCP69XtOnD9OVlpYw
XDjLH3cEtRjJOyDVhCo+WOz2vfBDhaFSVCNPV7DehdjnGnSq6ags05UDzqoAuaDp
tQQ1ew4QPw2T2Y+Ll0umxNGJ4kbMNqtPQmMGSsKayBhz4wFmU7UIjMhLyPAU6ggg
cE9wrLth5AQm5iFTiIX3KmNCYXefo4tUTfp/fCiYFRvbKvrFr0Eyujm1JFY4g0ib
LFpVR32dIc3OY0hoi5v4c4TlP9zNQFm2X8pXF5n3DRVteR32/xN/ZIlVwSFC+P9G
Ic+j1byH0tRN5Ge5PPAGq2zDZ0yUSzgAFrtp01m+53IPHvZxhWrO2wUZ/tBKQ3qY
CQ3QkXVGCyHFTC1MjbnP1TEG95LF1dmIfF5nVIZxXyE5fiDR9VG8ppIQYVkz5brz
6udaWDc2FOapCloeNo/zEybc3q4x3HCcyYEk/fmKhmIDk/XSK9GLo6JsOvPEo4cC
rP4dyLkgk+Pw3AiOD0oyVTG7M6U4YWijyR2SPIes86QEDU1bs7iciAa91CnK4ifd
wnizJxy+00ETqJe4232iwcUWaOtVoA3+V2xbHyAvbraMDtrNAKbvZ8cQCa9bVa6K
Czv8UDwstSYL+dX1h/IJ/5558oxcjdT91Bw9v+KbMBeRAuv+tfDCxxm6CwHe+CoR
0S7mbhvzNDRMJNCoOUj/10ra05VZoVLhASnBCy/598QPJ0UTzi7C+OlY3CEoRE8Q
/8a1tFMoy9Y/Fsypux+QiOto9tKW5YNQM2w6wVHsw6I3FJ3NJeWhk3dNrjBQiykT
HZ5Z+i7GxC/AL4+CBT0AlDe4xu+0toC8h6MBjbkpwqKOmkbOZCFz6j2YhwwKZQzx
1Y5opmSA0OQEGruuMqP8kVgIln23EmcJfxtNoGePECGkLQp4awr3boMlgZkp2xRT
jO8LSJrNhkL6nWqbP+pZ+fVPkvhaJAscXRXVi3/CBeuPo0f4rlD5lsvNPFyfg2D/
4lsDLAS79q1a3etzyLrs2BV4ejOqzwv44lhgx3m2//StIS3KZGLSZ6aXnNzJ8ofD
QLnWIqf4tLkoyA5tfKIs8uwspicc3uA3yuxBAhAkT8SFZcA1Sv/8YYbQLgu4LvLQ
MDfPP2UbEoLB+jUboyJ9lkpeJ1VwRLQJdoA4Hi0XJAe0lRRv/U0AXhJlhEKJ9RkT
tYq+m8auoaJBLxBckAo2+auA527wKaz8DGVddDTl4C7ScIMhCt46xKsxKAa6XpIX
uK+JsGo0ra/cBSwRlgmwhem7q3MA0wbV+MrRhiRBx+HD3Umyqtz07qoDNdPhDsiy
JjrX2eAiR5o1n7tiv9/sfO2+wl/tGJWGtjdW0isXPADqYMC04L5gyJbKJb7yKDRm
kMZ1X04uyTJkITCsp1Vrk+JlEHZ3QlPS0otdbLx8ItKG5yyKqzyDV+IXzN8W1YUD
mSqB4jIL8EXRTOoBUw4m19SsRNWIY6rekxTkjFOqJTlKF/d8b/cD2hr1ObdlkKlY
gM6p6bFvLndnWKD++CeglOYdRvsd6nLHozlA3ykvfco681N+0HM4DKmtKkU/CBjO
k0329/lJ97e+3vQGKpUHo8SZppoqZ8eiMgR8htVUn6bsrWHwXKTR7ZzmNCzpqy7N
EgC9Rn4sowYmTbKXdwMtVa7qe7OPMeCQ149HoGTdBWDgBXIGMw1swFSItdSI+jcS
7CEBlZAdBcnSM13LlOgbiP2fDcrfDFgzumtGdQPX30mTTWbyuOEUQncD7Vpye1+H
drQPdfZXfV9QpKBubut3HNE4ky5u5/l4gZtYO+VxfAoWKqV9pYU8L6ft+cFCsDVG
sxWIOlrWfUOlYyaNs4P87EKJoC+hDX2sQlHGUn2JYpC8Zu/sCUOs5VuBge23Nywq
pBLl+xUboVCRGv/rs2DDlRZaz2Wpq+zcb6DTHGZuzpxFZ7bjzgXPKp4gI3eRfE3J
AIS2Db9rCzcH3I+YV13coFSKP/FfKBszeCxkKkZG/mMpR/sliGBOBLr/jD26wsKW
OEtEeIoqlcvWNANoqj1+dC02AYAKPRX9W2saMq3hiK18XwK4NxyGr92Nud5Y+kdt
oVvULb0sKyskfWc17G+EG056q/uIMzWaptBkFX/z2NWVsd6CVC9EBOclK5k3RZSN
G+gDaWM5Ec3i9gjZ1lqA2bMnVSc/JXR2QTZ4R2yBRlbpOSpzMS0FSFaBuL7hHmX8
l+t9sbnAS/sLgONSKwIAlxmOv1/7bV/ZQD2EVnE+2a5h8+Fo4R8VSSROr54CNutH
+G7hY/2RnZTg1ZqPof2TDWKJ+0m/yX2k2nHJ/GNNefKTeaf32JcroiIRRqwRBvTX
JC10FducDtpjy/w48wJ7K5h96L0QPjswvseusRmmk16ceqTktGQ7W04WjVIjqvr3
9uBTidrt+w8H/oJpix/2i92yEoovSagGd8XcefPPxYYtYv1UMEafnka+H6y4/zQG
JMi6xjHpLVpsDBf9N+toRbt8THTFWtd/QtsdOkecviPPWMBPf5P2biTxtrgQYsla
oqbjTX3OBbxBL+M1R5CMw7DyFW2F7jI1nQnowHyOCQqB0K+njSeb+0c/04Y+I5NB
rrhNtzNdjzmiLSgZ0uuQw7S9Sz0AiMOvOx+H/zRSyk/GkasdebeKv4E8YMIpmk37
NAU2GMFbLD5qYHHoKJI7pGRUYU+hdYp8JYwmyziNdVDuXNt6opOEYOaxAzJn8Jtf
MPxE8VU5wwr8R5Fp23Uh+7wGI+KBesbM7YDPun5H6Iy0vMcHhWJxx6V4PQ6Ssx36
M+5/+xrt5hjktROFIifK4264Dg+f4y0RcSQSmBgL8eAFO21div03GR0in6+L1UH8
PuG1yot4Okm3HDuATRgEt438C0Nd9W43rwScMYWsJHJc886a53OqurwwYiDWgUu6
7TfsuYahwrCOj7QjWndGmWXdpATCbTF98DcUXw8VnmMQ3ASLE8cOl0oOav0OcU5t
e7ILQ4DRs9yzQpQzuNykhjeHnI6Wm0k4e5XE46cAr5H03Qn0YLhA60mhfQ68w8jn
2TC6IdJxaauGow+nVw8Im7TKfF44X3tpTx50eF67uZ4uViaYd69JksqSpVTBt5vN
sG0ZlbtSf6ijj0q0vGuGHZteynBGoOhKGSLOyZ5B+VhhpPYIW8x1Zc5qXoTx5jXM
dEXIY2iB1Lir5NwoQw9FLutKoUXjxPAFp38mJhUa8MZtORbHeCXncYH/IIcO1VHm
n+GvxAcy74HcQk0phLolSa4TPLuPQN8J1MAEYPl5pDPAcAm66e4GW3LMgveopn88
sd0yEz2ZP5bPo97BSYqu/5xdusrVqtui5HPdn2EjFLqzmB7aT98qYDFofpC6M2NF
nEPUjx8pOAjO59ujIsiZy8nPu327b4aysD+am0L2ZiCxAN0kYOxjCeo7ui5RvwDi
UXGLFLc/vpAcUtOrY0DZKBT93vLAlh6F7JG2QU+M9+e3Qc4CUJRaFoYDqr7v1DB1
K9ZuEFF/Ko0XX3d5apuH6pNHB7IQ9TLE2xwR+/awQKOiYWgtk8ImeJ2eCoc31PQ7
sIOScGEkpSRDf/33xr9iUBy5WBEr65/xgWrQ2uMsygscomtY95wnLVAtkpCpXq0V
OkJ7Hm6fqi3BiAGC8JTB4d89bjyV8uR118thS4kQsDgJYtGL3xt5rmaWW9B9WKGM
onVwtF4EQyZnLWuKx/4LON9U1FdAHsmM05TCZuhUlAlXL7+Vsj+5Qb5LXWYOZePr
yc12Og0nTKgEPwHQSD9FsgSX55gp9qa4V4BVXEKdQN46XJe1RGiQUDh2KPrhktH6
VF6xle1tDQGpyoa/uvTB5cfdENCrrCt5F3IjQFiGoRfTL5FYuy0hgZXrjSxXunkn
+odh6OCua058B6gr4IlmrSZYl4xaUA6a3N1bdcdt3CWDVcfW+uvndikf2igNsbJj
6FvpdkpFwY2PsKrmdC78u7Mt2QQtROWfaiAGTAsuxnZ/KVrhAU1lHKGm9KXqvzNl
yqXLyrYCcN3/azxxiqAxnHqewP7Syp9wYf1yw4lE1WNcCnPVm/bnr54A73uYmmIq
HuoiiG78OiqwdWc7f+72UrxFAJZaorHwvqJAzQ55Ooq4DcZr1qbP5Xi3L+eulX4Q
5MtJAZKbaFPPHNXg0hGtzrQon+Nb06dkbT0rYXM0PTjg/c49je8Ahr/nD7Frp53c
O3KGDyYBaD1EfBxVSL1kw6OShJMWH7inQi8Bj+88ts3JNDxkiH7T0PEdmW1FLrEL
h0sMa9GuKjVORwLiIxdqFCfjcKvq2iMTqz7twWmi83gVgnDB/GE1ETfApgESImIO
70Sf8IyCmT12txFpQM1WySnQLenHHhfv5gpnTxASugpoAxPLX3Q/Ghlnxj2IN0a+
dPQkGXTNqbwYbQPv2SXJ45x07kc1PZuYQ9IT6IrIQKONqeN/fqFm0jGzpPOBLTrO
7TuOZN4hAHE6Qa3bSa00OH5khL504SSYbJ+oQMXNIDSbLUdDQh0iqqYQ+Yp8NWTe
uzkZyMFOhAv5fJoyGqooD8UVKohs512kMQIni69AchtTVGFikN0f+8ZUc00yYOd6
nQFtOzB9bHewztB/gOUTg4braXxtchNZZevVbRmMUmtDHCowELXKE8QUuLfZiqoY
gNcQAWM2bd6C0pS5seSAK7/xIYA8SeSV/BMBG/9ZTatat7siDSUqgb+TEvvFQLsE
ED9NrDN4pnNrdb/letj+BFf/YPH8DkjfB7Wh0ToXbGlHuPiyXkN0MFhO4cjpBXxq
4dRJolNSAXvrQwU/cFQ8hS3h+OAa6Ey1X7iHtXPsCioLchteN41Ph3EexwRO1pa8
EjLwqrDnTFoWlaoE6W6Jv4VLV15oYMf8/ou7eF9ycr5tPr0GHKvXN0Emn3/gz8ub
Pj/ecNnszuDu6gOXc8f3plJcUPKE3ORykwOIkrrZTvmCujhyx8E+xvR1YxfKFc6K
9XFhjI21yRM5oJ+Of6qZUjS2THY9abXU9XoOHUY47Oqf46c4URjIz3LU+HjY8fAG
7ohQnipKKj5k+kG4+mOKYieDtdnEXIiKFgKZVLZ6ce/P2o4uXZM1sqvZQj/W1WIg
e89SGamOjLGAqxM+m9h9naeDIp4w4Td/O+JnXDdb3Ha0QtuqoCaHbhq7KUZasKsy
WpgTH06PHCl5G6zwjTTQNO7cvmK7A/JIPB3l/l+63p8fyBqfk47J2XaEjoCv8j1a
P7uNXEq9YTCENXR7w+erEJhwTJZbC0Q1nLZ5Z6061bjgeMQm10GAte6m0hptz7Y9
JcICPwbCYc/tdpByETZ2hSZqticfW+OHgFZXbV0yn/fsaSKkigPgvQHJcw7D53CJ
qE04OCV2d3DrX09Ohjq4s2QRESFfx6orGWEUuHGILsPUEmCjWHAkTZTg4rrvVRWP
9f6jJiorO8/OEd8HnXOtRF2K28XjuqO2i6DEFH++/rtPCwzkhI9h6+7QPD0VSEWs
wr2vqwb7DreMtXL4/Dpj3X4d8d+zUWWGu88vEBl9vtgb567W4JVV49zeU6zOwS1Z
XBIzxo+wkZFyi8J0KVeHN8ce6otw88iA96IhsL9urcpfLaX8/9eZCrgeOt3VMlSs
gu1mryQwSpYQbqOEI0OIcgg6XmSKWZcjL64+LZ8CbX9O9slY0gz6BnhSe+SP751u
6sUYUUNnq9+qWfqB3ttC3El4YNS1/mlST/Uus1qsH9kfPZCEJJsMgb5WtIj2DW8d
YAZwChkgAOlPcOyV6DDiYBM5hIa9A/0skF9ca9AyP9Gi7GUv13LTvVltn8kh0w9i
kD0g+SGMbVwoiRGSGrvUmyFeaslJdAOBy17tNk0TfFnp06QJOft57eaJp11pvB1z
EYgU56S4sWDtA1d0MQtHGoNKv86u6LP7Une2V7ptEBvzeDLW/X4jzk/TqM3rZcmW
ZLFnyuwbt36biEAiN8eP3wrHqkd0iXyLKYVcQf1HU5tRfVGl14Yacl3InNPPn3mp
MbIaNKnSsCdfwOWFRKfNhljCjZCmbn8lt90vHqMrSh2osOdNme3RHnUBc+UpWQyC
eji2KobqZc5awNlc7nGgFS26O9OgpebmKT737DDd6h5ixzgxE6FX6X8g15iZnjZj
44ez3GksNF6t4UtF6xic2PmSHTzjV25ghSKlXXqNfQyNzbLxpwNG3mglRtcHNdh3
Um7Ur7W1uDe0nv8Xie8NVOOQ9k90hZ6VosSevPQwCW1Mou2jBSBCySCgdaO4FjMl
ijV5F3eFMdaA4/zBrVmycJlGeV2XRTVbdl0uoi0mOETM7ukYA8Zu09Rb/v4Ylfxy
zvfiUsGCWDeoLYMYi1h7gDbCEyEdoPHIfoOSZOBkyuIW3KiKWKGv95YE9cVKax4F
3ZXIJFx/zVOeaQlQQ2W01D+1JR+wkdRx0jCS7b9u7VGU2O6WxRlONH8JJYu96S9p
Qa+nqtST2gL4MTyh7JvJlQWU7vk5ZWn9Fi8AcN+dWtB1DFL2tk9wUCgqtFAHhPPG
81jmmtcfvPqOzWkYGWmSfw57Zbq19GsgJfv0sbmM3O/5osXBw6ZR1W/FLaihlOAc
aIXVbGSopPjRYKZjVDXMA6tt/c9kYUB6B8eVn3F+pxxBgJ55XpWotsOSiG+W53g2
UWbfXgH5KKrXxy9tRaq4nHcdwdA1h7FnQwmnjqx675AHLgXLtD+RdEdWByj7BLjG
JU1HiWyW7ZlLfjoLuYQQmRM2fzAxtDL4h4vrjbhPqtxoEX38JglwW7ewXLjD93VB
8kJv4eoz52vvZpqwpknjZxICXnHpBB9OQ8VsbXzZfd0n81z3stmJTtZz7bMhRGGO
Kd5PjFJNMh9hK1hvwq5kj50DiJmt9KA4iDeH8AK5HZIha+5Lfjfllb/TuhlmcCa4
e3IqHgthu4DKoh4lShsUjS9VgR0rRNFTeOCM6cdcXNRlLvM2MLPkNdS1ciepNOA2
S8U/yRojxHftG/jeauy8kD8+yy9gPG0Oib/Oi76uorn/cIPSf7Kpw6615s4rC3xj
Onr/gHAddq7EIJtFU/NBa5YkXpXy6fQQhshNEsEdPbaTiDEUT69LSxx5TZlkQvVQ
7f2Lpidzl5TtZ8PL0Qn0T4pdoWmK4E2pCdFu5eY1l8+cRmWYiQF+IpLPjkKKYDFv
qC+LYI7fhx66mM9nQGku9n2JKd9ztsL0t+hF58FIF9Apj7x2CKwYDOFA1z9Gd9Wg
Efk6vEvXvzsfhXsrOQvTyQCi6pLt0QBp5HVORWyaiR18mW2PS5CsdlnZP3hgYPPe
Jw81fvZE492Om9TfQHG58i4RY9PQt+tcJ6lO7lx07hgkQz5sl/KHhBRgX0YKWiQB
6BRJPR9i6ODfdDlPFu7ctjEecA+a98d9c8YF6FvSpuTl9XMrg432zETiPILzzy1b
xn1Q5iBfTji5U4GwE3z55qK7ksL9nzHVAQ5g5BTG2VLeN3uUQI7KRWUwrRTWBqkE
RYzH74zuT0AiSfpZkgqbo2IxutBtThj3NzXXhwhCcmdLT4IfhCdkiZqbWCnolGdY
cAlT9enEsvZu8+W5UERzRCYUS1oZnuAJ75KASNgnG5PDV2VgNF0CyxObuHOQmXdf
3Yrxe3JUyS4WB2QIiSsGXG31W9IzGf7VehU60z62s/L92i1bDB6kUBN09DYpoDIM
UUq0TbrSavwqWabrEbGUpSGTVODyZnPCevU2kgeT/3gIyfbEVddEWGh1bz90EQSa
InhHqTtKDQ4cJkK8fvCpSSkQaHJfjqMI3Qfux8oCHfxHxvPi5ACazk1RrA3AAQDa
f8f8dnOWGjbWE/n2TiyUmJKBAb+T6caI+1NjwDD7bzXSoWMIEzvA9U3AOBhQ8NAv
1RcWmOGUwFzFuCiLKJzNbfmgl2yO+tD+fFWq8w1V7jliBbEar96GRiX2F4bMM53H
5pefRXVCqInGLNpbV+DGCpzQQktP7QKpZLNUapAbBfMM+xM7KHTaEs4XJM2Z9wXY
WbvQx9CPE3Hidmke9wv92Ef4Fcwq+BbOEWG1ElCFOzz9IUcCai6UWMU5fORGaiXn
VamgTtPpfeyhgXjJU+a+S/H2Z6m+rsedkCKP7qtp7p10bG3zr5EQkNYht+WWNoyY
pcphMKvzL/FkNKwUHCZBDqQ2OPWpB+5vCQwyjLwILfkM45H20q17Mh527kgoTKhi
UZlXut2Kw2pXyPYx7WV7DjXAB0BsbuHtAF2xCt+NE9z3hTJn5e3UL8hbaEznB8h3
qZVf20xbNLfXuo2duJPXDJGKDP3bVAhY1Fqwn3m45hRNklJeSHzR2Y2GeSXj4QHM
422WTozvss8BFQQgiIO7Il7KO5thc2favmKRsVhJDehwJJw8nrKpzho/j4Mbfgju
DC89ampcb57gQ69VZYlKu23zW5J4bIg31R8zzidypxtuA3JA9u+gQ0+TlffzeGik
zEE4oruxVa/B5dvF0YPuy/wGL07QqK+ZNnIGTy09pBy3LYNUON/RcBcHzx+rcZsB
+Yv7oNRjwRIV7pHcTMBvbzxhaiAFl7bNufbVq0AH6ktVNn16/n+FDR6evN0XX5wX
aRSXALqcxxIWXmH5N262IQp9CB94ZIxPzJj0IxqJ38tzbIw4SlATfZtC3UvZZ90S
l1C6EiaiWIvQo/fqX6GN6y0fCDdVfrj6Nc8kTSjUng4jlUAZtieWiO/oSCR6G1Ma
O7PvX7o69QDYqHMFFg/uS25XjaHm4nfUdfN+uK0XILxYlp4eCdFGDwrtjnlV6RjZ
tP6DQ0sdMjBo+hLElGaHwhUqSGK2gpAYeVibQEf3QcpRPiQ/Arh3tc2PO65jgFrW
nvE5LKh0sV/DE1IG50LqiXecTDqJGkTWMX5580dxxlQwiUbs44/YS0MglqqmA/5Z
Bg6JMMoGYO99dDmOE53ex3jk7VbS63NE7r9yZ1G6fMocuDzWpQvBza0aqYLU8u0x
bbNcQgn9gdPPnKQd65DuvSF+s2UtuZYCAm5XuV30GH0r+Zf/ok5J718TeAyaOuMN
BrZlSpNdETJH7S7/+928rfH1m26ZIUx5kGnpRgcisQGx9s0r5oepSJtQFmxm2oWI
638DkyA54hifAEiUSIv4MVonYsWTtZuebDQXYC4Y6CnFSxfBJTMjvZWDHjbqHWAW
jGEQdJz0ZYal2UxnmuErS6PM21JbkyCqi7cyzyGFx2kWfGAWYa6IOBARNG1PHYqM
3xwiz5gbe/ZT2RlaxSBr5rmZ+0tlcQB3RH/HShzgQDRjURHYDEqJVojCOnAau4fS
Ob4Zno4H89iH7sCeUR/vtWowUokIHXiFRM09CuQp815C6mtz5YILptvUKUiKxTX6
4MH/gFCQ3n4mxFo1gzHjuYih/PgiZ2u6ycLFVNtX6Fo4i/uX1kSK/JgaNLj8+pzC
kY4tUU062JLIGp0LCNnNEqDGCdLR0FZTAySSWe95YYGneBkTDUwlRyC+7yYYSHMz
AfsFMtg524v6kKYHjWTO7R/7r5mZeYHUu7g4ZuDl3/e+aHpfx8ueQmh4EbZK0ExZ
bBvDzozbozS2WlXSL7cCJGunt9HIy8gqKifz5LwQWL4nkIbcCR+/d2utz2Yt3Yru
Lv2y1uyo6YN4fsKk5RyxTfxgXbmctOM4Ay5XRLPBx5vgWRPfNVoPKv0C2VtMSKVH
UETSpKfNm9A/hhrJPXhcjx+BMgHzPLNbbsaaDV5BaWhgB24l728e3tLe7Ofag0q+
LQX8j0etON3DeYSdVeyqI38tlDOpKMju4hLbwGZ3ud6Q/YCEyNThlIswAyf0hs9E
7kGTXHtfj9R1vh5WtXYyrxQYp2ixD+LDLWfkFrE2y3o8bOtSEPOqBFN/4UsSWCVd
dk8pTX6EIdDXMN9XT69YTahla5bIbrWxU1ybfI613SAaPquxWMSpYWgAoBa0SXIX
R67Tb5upJvOEaFsqFssZfJY/HjnpmfXsPGrh0UC60e580KnAz4NSMnD1VXZRykty
MNz/Qa95c4+lMXu0Vbw5sgOWUvFRaDJGdYKAzLfCxZ62dMuAN8rnTAY/t4Mb30dj
/t8g34yrYhJCeRAceLLruulPEkP/D64dlvq5Lc77KT/vfDwRJiIKsT5MWHOuiUVB
p+rFNcejSEbv+qqiQj1gI92wFfIY9mQVmLSMk8fC4HX1lr7WJ40JDrtnpwfWVTrH
FjIypCxvSaPqqTYrDFU5I8jB/kpAP2mbZxGMD73/Qtx/1THUfV1rHoEZ3+R9EgM3
TrFpmy60LcIdeUtnqGf6278Zq1VobxUacq2qwAJ6iqZOXebOD7ixfpzgZlfff0Fn
04yN3UT+NotWA1eA/scceyvivNaKgXQ0pnloeCUgnfKum/nWADeV34N0zkZBTY9O
WiJuVVGFPk/qNb2BN5FHhvxfzNY2Hu9mve60OF77xt/FueG+YGdek7b34vDssGl8
uZ1M+u3ZpLS6/fFpVCyyOYQguJhfVenpbZ/JLrKcxiXC1rLgMAjHI7xM2AFmED43
g9OpP3I6GEQ0xnWIBR70zRwlxPqIF45e+/7phxYMfyX8+Sricmop1RyleRDzHAFk
UeDk795EjfZkXQRzko2kyJS9lb8oLKgiF9teI1UDCHQEUYZWQC6EpQPCCTNJt+6M
Nl1icpSTtXHrffIkE0tJU6wBMxken5ExDaUsamJXIOP7BtO0rCwFl0nR42GxBnCS
QDz9r9jBSysEQQUCmXWHXaWouG5mLltHshSNRdDEodcx+7APOaz0hScVjx3ZtFIy
YyK/k27jhIcj5DSNOaX4s7SGMV0eSY2NdD6RdFEF+3PZmD2Rc7WaUlqM/kFOBEyv
lRTZv/WEF7rXFdwzOLIEnfFNVIFxWeneFmt1NuiISrD6XxvGnEO37ezxXUqgWklr
MuXKW8IRad7sQiz4rjl7bOfJdqKFQ92MOd3l964S5SYJMKSVwbzOJKuaatamvzuj
K8e316PzkSAj3/JrgL9BV0TbQu8jCJvG87VIqbCDzAmWB7Yys3U1uDfjnpWZkxHr
GcI886WCcosoJ/moe6DRuSnt/zekro95EcX12VHTRZoxzVGnER1e4+q/v7ygB6a9
JetQ3UllkZDFBAlPNDJ/TwJdo7Aw5q21oKjSqkhyrZ6mh0Xgz+9FR6owD1w62h89
HWDHv+7GHj931uhHM1V1C9zEFJjoKbrnWgMJ3G4y6ZyseLF2TcOOsCVOzA/QZRuU
BE3WtPd1dj0WvVUr0XOzEpmFAl/5PJoeHrKzuF7HFMRkujOf5mMpF1L6Hqui2KUZ
0T3ITxyZJZC9TEHN1nel1NikeMkkY/6BWWNLKIp/cRce2US4Ns2MBdj9u+wOgMp3
R2dACt7mBS2EzZe5R7VsiBkRpnk41QPQRl0sDtfYLhmHoHvZQGWQu9khNA/0bipl
FeJRJCRIjBmotljwMLSY5kMKFSPgQQPlCdOHsD8pEPD9V5aGo5tKN0Da/IfFMUWc
utcFGdWo5Jgy8ZRQ4HeUeht0WfepRJDgpkvbFhAmVX36W1nmz0tvSMvL5Tqley6m
bjT0ZTxZgd6otCdNDfz5q56TWPsa/N7013qVAA09xs8Vz+5U+BwACn1utU3Pd5iI
qnRhdhFryUa/39FporSt+gus+PabM4uY+rEwVqk33TOVHHnUlYvJBmRXQ2zcGQGF
Ba8abP2AvHKv6rDCJBeC8Xdxav5jXc4KLZ6sH0YlIMuyiJgn/Yk2VBHi70C7TVmJ
Gy3lzTugb6j4Nch/d7pZ73uuKIOz0rxzrBjqPzoV9y6L1sKNezLobOLc+17X0d1m
NcFSES0LD+j2Gh13+2orKPNVBjdlAaap0pSU9tlGglq81dPYhaqxu2D+wCCRKXaT
K1HAg2w5KxjzPl0O15NWGl2CgKyAMkIB1ZzcVw8vYBtu9LFsCooFXRlzpmaS2VF0
/mk8zYEnijdS28EvsBDJRecqskyNh/HH2/VOuXMlbUALBsZ1yLRwRo3XKV5rAQVf
PmwW/urZXgZdij9D0LanoH9boxqXwDHs0hhiRwS0sCO3zSvT/1KtarBeoUm6T2a+
lF8zVvlbuu8YKHMUmb++xY+CCBa+mL0Hwvu1pr3kpj6reJXeL9lnVKL0mljtlDRD
S5+7FD/OH5yu+98DWfMjeRbYvcDChq998u1W0+Bbq1LZgJc7XGL5Rhhg/s06OFB9
WClOMltoYVLiA6DRZqR3ffvdLfLDdZlAOS1733BySU9k0v0kp+Ki8Usf/RDsHA5g
WmHbQRnb4L3+0PM1RW7mCEnzP3QUKQdC4gIK1pVve2GN5VdqfG109wr4UzOMEb8c
wN2wmR/4TM0i+6P1KmIBujKof3wfKPaCxWf1M+SyZuY7bPZge2mLO8gq6Zkhxebx
iimNKNGG+oa5HeYlvKnIfBaXnoVSaDSNw1TWZ1qbOAwPIYG9oPElPxGk6coBUzmW
lh5qQmp1rPGn+snDTF+/lSzlrqC/hYsr3wVZxa3IU5cLvDq6MSnczhFm5GW40++i
IEM7OiurmHutZtCm82rWQ6BoYYe+hm4RQKpi4KtOhEpcMzVwE+1oTAAIAnqVLfzK
IBhLARUAcIbEWmH5x5ID8yziybjxX9RbzbRfn4lbjEK6UwcX9DVc5tqTjbHeTrJT
KbdkP+9+D8gP0Gdl8uVgzZnT0LBMms3ux1LNh2Cqj/blOKd2xCe0fj1OcSGVjzfH
rZIEe8i4D8P5lRXmOIVbQ9Yl7BZklYtb0XMBTXQBbEtOKirzEMM9ZUDpt7e0sibB
rar1FtEU2k2XHzPZhxGBI+yUvZpw/bBJolsNbQpugHBudXrMLItDTJwXXmE3Ywlw
ulxmkkxV4EitGD9SdxgUe2Z9EErlqAS6km9CamlbYIMfxp9tlWGSfSN3wYdMCnKC
xLva/S2eEq1c6SZwySJLI/n3lUzNA2RWG5CqL8m/0+V1Vc/idFE823/GUeBBE7Ud
9NwpOEZpAKKKVvKp/vz3Np4clw2vrsd67OB9ehrNOxRd2rF+GiA6s3fNIA01t70E
tqEVOvw3BeRAxeCv9Ct2A5DP6YZ4Lqagd4eLS6G+iKVDY2UwEVB038mCdxjL2EXC
fJPt17O3UNfYIAPvqLBwTAA0WsXSN3mpgOR3JYnd2A8nYChnBWOtSTeqhDMNWi4M
E6pgvmNuJ8vNumPciF96OLCEXglCKR/yCeyhPqAN6pHh74IkHlDec5W5/GaYjQZF
x84TMkgWgFdqpmJWhKCSZVDZNHavJGDsAaDAMSZjYIokinBBfi+dlcAf+NH1w3iA
MnzE1xFuCJZY3zPozWZNblxFOuAdgcigbxPbP7+CE0AqAU8SsqNRDY8+1Z7PDCrR
/wLp3ifGpHd2XHQPgdFDQOc8HoTbTr4G+aJ7PPftVBSZSkijOk9t5sWHr1uvckF5
a2+8H/rp33PyTjxrfBY2F55lf3Jmf8XQ0FyRtfwJOuhHz7uAmBRTnBjcrtlxCdOc
HNjsMD5IKLaYGyZgoAGoXN5AMq0M31tfHYEB7UGuLNr8wbrxHsk8xfFXF4t3SSRb
5YT2WMniYSI3OOy4QzI7shjyo57dkiNPuJ1KrhekXZr5pSevcgQGeldN6zuOA/5M
6gXTnR9Q1EssCrjueEhjm5QbjJZwgq+w1b1flhkSqFytngQpVIGctH0VEvGaVPVo
2drVgjM1M2o8hrwnTo28DyLTBQNGlwJqHHyL0a/HC8XOiOUPYw42Gd3ouwC09Dk6
hw25UmaraL9Fv4H4kDVyEInvpf8RGuXYy5ZhV0L5acCynoJeT130VJMkMI3Woggs
fbEFuq18rSGdCjHcbKXQsR6dnfLwx1VbAs6CQFg1VOiZDthos9yjLopCeiGP4huq
9cP+eDNSX58EnC2dt87ErEWnce6diGilFqnoRsHtcwnoA1aY2IMzzMQbYmCZmhlh
EYV/kAXFtipgiCwMkdj6ZdEobH8jl8qIP8cNsKK3eyNlTEVmvvFHiFUoGf/PTm67
mZV508ItVDRXyyml6uPGkf80wnJ8YPAGi+n/9cSH0YG776+kcwEbgszJwzH3orKH
ci4LrHpvRcazk+5xHqQN4WUy2Fqlnwkb6xLBV/f/FJmMP6kTrgr/MuzbXP/LMncd
wh4mRPuQ+eeC3pNFBu7KbjvqBh6I4NLC2xhaubrTBCzZsZJ/QdVNbtnGEgbWKGdp
yaOGQfVuDvodxeBQfPLRZptQk4kftL89wpQbAOcIHHWvS09k6qjSlCxLRMejcP/9
aaLCIAIXvdJyxFyBjemjOgdEXtFB49yxEpxJVbwM45PJC4TcY9zJ8JpeR1BFDYXI
n+H63hjvwU+q/ugz/NccXPQv/71IYNcG1vAtjAxjtS7w45sG/PHmg5o04ahtrWK/
VXVf1UNeXmdcOVa3OlPVdONiUVXNGSJ+CthKi9clBh6I3A2TntWcHauU0W0DWH1D
8RbRDr0KtYu/rJHkuaEkBEXzmSBLtwVarLWifRaFLTJq1sPlg6Dc2lC4PAfe2U20
Y4ZhDOngVK7TNMH1X4hEsBkOSgPbLsWnSZzQgy0w0ahyR8N1evp6WgzkZvYDaOQG
YywhZztfX497sfBNIW0KLRiS9ZJ4cBdrLPJrtsR8BCS7Cvsb5WPkeiq+lWao8eae
N+eXRnjgX69yDqGxDm89CC82Hs+QrAX1m8N6bZ47McXhYyqT7917DoWGq0t/y6we
kMu7inuSPoVEHTNjo7wV1BokGPY/xbq0FoH4IekdpNcgZFZK7LYoDb7CuOmh5egx
nxjSdOX3o8lvq0mT8PQAuaPT3X//3xVm8m3WQH6Dfr2JKmT4TKRDxCilNH7eIAul
ZTrmZTnbdeaViNOIsN/vWnyqYVKSuZVDajWohIe/mQe9qMPPzr2Z/GzERhsY5hYl
OdA8/DoPGfH3NJXpQ7mGBJ6eotWcgUaM7QuLneQa1z1Jn2PhAJG0OLsk+XIUHr7o
jE25aIVvzMa4NlezFUS7S9jpTuouco5d1Xfsqvux3QXpk6yr6p98BqSjx5rhq0RE
JcnCi6o4kIODE8eEB7RWleKtf/JN2zmd6g0T3BQLnR4ZiTCElJ5fYlenwuC/Ofki
62uz/lKkAy658QVeR7WNP7Dg1CVHrVxADoa0sUzVrrVhlDTKEq0Cz4vubLAN+WEx
3lDZAFJ7oRzmmXc6hBEqFbPLKQym+4nfYsAA6D6k+/W/q9llJJZmreX+9E5tkqla
zIC+wUYt+TNZcZbf1DpqzD4QEI74r+XRH8qImjmIxQPpu3edIVSxvn0LPgHulT4s
u9Afuf7w8L4/UAReVy5MWqEWbWkNkzy/MiUk3r0BF3dXwvFPkqLoGpVk3+jUJnuh
7MmUbGCnj0CESTfa2VezKktTK5ShOMoafBMna7oQnBoYs7d/4/ZLBDBNP+jLx0Jx
RToFcyIeDRzvVlfgLASrSDGIFb0jWij14DSRek2EC6OLKk4YDlHhGdIXpnwwvms0
MZMr37H3ahZZ/vsP7Xt8ThtUPz5gFTbncg37nZeqNCuNPxRop/oCM4Pbm7QrIHFN
D4fcnMEUz/CUYEPPN3Pp7Q4jx5sQSaQIkWC3hdgMZ3a2MvD9xpBMLAPbKfSiIqA2
TC6LQsv/eyMlD7Oka381Brwp4HfFh7sBns0ZZvoxdvsnexAqmgM6MXcGPN9/jd5C
H5DboWTdmLA6D77jPE9MV7IbOQjlj4Vsj7yxmc6CvaIkaS2Tr3Pr9PTA0KGD5Zxh
2Zd9eWWIS7O4c5oh72UUtMvS7ZKxZC3QCw+I4mD/plw+2bBUlWtos5UXo49b7IMS
nvFiaIHifHOsjeUVggoNqSlFaPz5aWSnclIsbcsK2y00vgwP3rUNnyQ9kMrn/AtC
pRQV0Lr3QBXiZDr+J8N2nxl07ALaYWr7OMPGQaxdscY3EWC3fDDcRmtgU5hOkPUY
FhkQIvOAoTkTRTHzpDYbmV1s8x6HweaIQt0clJ7FQePEHN6LiLG+ad5VUENWbPSw
BZYeAuLUWZu+27el/XUNNT6ul7di7ZbpTSgOKchfazUS7oZW/lkpSoioZsCPkgNW
s1bOU825NAuKdnRGoM381aEjZ/exf5hQxdzn52OejqM9ApY3faGcGhdMh+MLWJRS
628x43dOUbhRWR3HJJYbWMDsVlRgwMHUW6Vzo3DrOpQvlXSznlosRnJqnkzChpKW
JujNJo/LSzRQbvUbRplSIwlzoIK0WpF6SQPD1cNBO59WIeCXjDY4MdwxGgIX0BWb
1cfEccimFRmYH/07oW3Oocwyc+VQSWPWDuX6Pob/6kpiJ6eQI+OM2Q5HFETrQDlk
G0DX4em+WMoY/0Jd3ohWSaOVpNHwz+L2k3HbcaJ7c5O8vRQMEk5027M0xaaxP29h
noTW/3U8UywvAAe7WyzDROEpvUVSU0nUXVXlcT2uRpCIaiLcC64GmCbnMZEcGE1P
rYNAhLo1MbJSl4R1zpeLfxaFyWW7spxFbLPoSx3MgLqz+V7DqwajR3+VYb3ZwOF2
VlIsTs9gTwWBl7fmzAqt6rF3AJoU6qjgYIkAknai7fC7ZGjUkRjglGAjJmDkVZ5M
ksSPVpJqPUrbPKPy++ghY4ba/jFGz2lTVaRjrcuNffNXoP3iEsZ4v2zUyGbrsSj8
NPsnvw020FND0qF54SuHQg6qibnFd65+5lhAErrNJXiY5llnJGKyDCG0yLYjlGtv
52lyBDmz44UPpcXFEmKlTHAM20eTCL1pFuc5xsXhVntVM5tcL3lOdHyB+StXMX6n
A1ofRsfzw9nprprxnE97GA2MkzZci3uV54IqhvhNeyW0kTewKayHiFwRM2cFUosO
KXNsIVVQ6rvoDsq2hA01Y8gT5sYv65AaG/OKMtOBtcEsTcoeakDbFKcBfTNbfSyx
v1EIo3M3ImrAqfKwvO0Uv4xeitP6Tx6bWFsdlTNC7I3358M+NFLGYbr5+QE2BHF1
Sq8amzGYJMULWbmx49z6Oktw5gmI8v4jyspnAtauDH5+JRv16UwsP54+UM6SJwwa
SYRKCV+pM6Ly+AnjBawuJ8AGWZL8jyJNmvjFvuxJe2U1IZGzaoXKsY+ewDoF1nVM
kbnnjV9njsX/TuNnnM6ywGW8eKXH5Tw5vNsulhb4ZLNHICjGWIAtME0r4BQsANOn
Cm71O1wgmGtPVlnVpuf3KZoIE0I3AyuBBcjCOvpRqBELo8cQgmLdo53lvKAA1H+2
COi1Bs/vNfk0b9agEq+Jjlz0Bi0PeND9DMYLJxujKAVfhu6a0oVFgcaXAIJpf1X7
XmzDq5+BReEOCj9mUDDdsTJRFFd9LZ6LtQaPyFpaHZPK6Pjsuf1Gku+OmOgJSxXF
O39fLDUUuKbrBLyWaDTbZTarxIEyqo3WV9pGgDWVfDk1BW64QcMrlJiLSRegjihd
TWVU657tSJgQyuw5lFha8Tp0+1zH8GffVb3eIpXdR7i2rVnoMbRnN3lA0qWOVVDZ
py/bVVptNyrfaPBP4Mo0nOKNYzxDp1n1FsdDk5vZbK+I4MYEYN2YBuJ80hFrl0mQ
KtFCjPdEpr9zxPLLNgm49jgy72IQyn1AXquzTFlf5MnlaQa2MlyoXK+hWsVOsiCQ
aOeRo/1e5C9DBt28VunwSSVFySRtjUyHwwECp/vwNZ13qau/yJfCT7bfo6pnsvI8
pL78NK0iZEHBMgc2w043pwCYC0zGQpTWTmQ5L+KO6VIhV3AifopCT+DLhAjILyeZ
VW630+G8eJtmddTkT8dqJVU6byqMuq8cKIYas8je8SwVMLW+SeLrHif4kVLajYOG
bYll4E16xYGn09e7tgZt5tFIwahaNBql+oPkM+nLWpr+nkdmK284qtY6qEm1MaQU
EMsNS7iVnGXpdVfi7p0ETU+2yqcA4tT/5vcI/6EAEYA4xPMoIuV74oEeIORN1BRL
kqkoPxfOfeZN6jpXDem9Fjh81LHJGQ/YvNCa409wySEmIlUoBoyOjNdbroUWD89z
/9hbJkv2pwCT85gfSCIgPJmytBPdxtjc5O1pd/3+9PjpTz/HPToIf9VOQDUMWSDW
pa9m80pbdt8rKZYXajrLXHw66nBiSe4MhVDFbyy8Q0CKEDzS+qMVaVB62fvekUC+
e+bW/u1moY0c7I+2GRUmAJ3HQuIEBiVlEK+S6EhMIu4uJyzRHb5mZ/FoWDG0CX0i
xORMkoUXvq/e9J/cfp53cNkr9FBtayrdKub6UYiwiGfv3i/FzKCF3b46L94XOpCY
m5eyYdHhUl/cXfGF/EgkmO9mL5xra9FtxmQR47ORHjF5OqmuL3gfPDoyWqBCa8HI
ziPI1OuDzayoeHq2duQqtXcnDaEO+0f5RZbxtBpMXXes8hang3HEsmuDT1TC+wcW
bdFFzlg0dwX0JbhSjmr64vKvq+F6s9cx+HN2JzTqxWN74lkVze08GjrBkDRq7vyD
jb7BTAnEnobP2vZMXLXV5OiPIG96FTW91Ka72pqe8xvAM7bEsjCmsZWpSuCoNHfq
Z47Cd1v8J48PH4cRSuXSWme99iT4QTaxTEt+aaz+n6LrDmgEo2qhk6/hBK++VKLV
40J+cTzhXtzgmskECEF/3exIw6tK27e+NP0lYUvYbH7MZtAMKc3fnr/ElfdmAJXQ
smx/335/VOIj+xJ+A/UG2+2e9BTdQDbeStWLjnBWvkgZLJFJf1XyzqvJ31lv7GQ4
+11Y7k9U66riKQ/VnXt+ygqQl6MQ0QaX0BsO55aGL+MxviIdl9ZF5duJqFQNAdaU
4qexdXiK9SdaE9sIQ/4EC/rBSsNo3PVaR7bRgLzAyppkPZ/kizo+tU7PxP89fIkc
+V/WA2VzSNRO7crCcSUhrmgYCGlg5+xVtVNNq0eTjRsSPJjyJAerJRFbwnrfD5rg
sm7JASGNU0yvqU2fwPymxro87q201XzfNj4Y+vu5InASJn3BS/AhDMldfLhcN6MD
NB0eTCblrE8WNR96tMZh4NdsbZ9qqV6C24J9ujgt+8zxhCSeXQL/+OIMDRXIf3Ov
ZaVyJh7hR6Hj+Ma4XE+U92z7ow5q5R77UwufxAhzXefRYRaz5u47sQo4HI/C1q2d
LDbwiOiEDqvRnUYdCWu/JiMEh8BQwQ7jeCHkr7GduFZJUf+2xOLPoHdUWOWDwtdq
BYg37TfpZ29F83i0cIJQVcj9Xa3nmtyFmTfjRKM2TMqF7nYxn96byXFyeAKdsdhW
Lyhwr1nfOuO2lZOG4nlfiFD/WI/Idty6rOESJZvB1aUbLd8mdPRaOGbzGMtW7TfF
mPVvLAF76Iv3eSianNN6PIpM8wB/4sK2Mh8GeLg5Rcq8JY5FqR+gUrwWhHRGlTNk
9+fY9V28A3CdV520BeEZXIRBkn6N5QIcuoMVBZm6cbA2iaA3sGREQalxDovi5KNg
zSKwfn4oLlYNQXLZiBRccP26Dbimk2o2ROB+1jOquRHFGop9U1P7U2fennTYmaYQ
uPMr/rOrFYMvclbv8dOte0l3zVQkpC4j9O0hRhcUtvVjidIX0tK7c6lLibtlvTww
b4ke5Itmil+LfHls9w45Xi0/XHMQokYoOkMKzlDe83M691QdAa1+P1UrtOUL/9xF
I2tiAZS1irJbBAMMRo7CTe0y9PH2/WPYC7jtGH4t2ZrCcKAh+feLVum5FIq41sBV
nXs57Z3inBUyTze+zPH9LlcahNGiaplWkE/iVscf9h/ZC/UdM+VTpEftMHt517ma
5pycqmwEF5GeN5XXSNyyBivlvqAyb/MIbDE6tYdgJJeILlwqm61oTlKQIdVxMls7
dnlTuUdlpxSwqMOVIuLrmsE4LvQhOTuBaxHdmMc8QOzXNMFL6ZournowBxdMgzaG
jGGe4p3ILMdZgyT/Q+OGkfb6pexXSYbIGsCUitOOecjL5YSXQN8YTF1z0kDs1vgA
Hceya4rilO0UHjq6iEL5tfNn0uLDcihFvQb0TFAhw6Xldu3hQEKWIL/m5//fTHI1
ZTmbMQTRAFiH5+d0RX1qef/HQNatMkJgy0Gso7NJwIeDuJ3XkKAEQL+RLSEXaizl
CBeUaMJusre/uEVUT157lPViapVeMdpwK+QN7DGM1XZD+h8lLOY+Gq7osdq2FCLV
kw+Nbhle0IvKE1rc6slvcR+BQsH71oT923KZQierxL+5qX8DiTV294tgx9HI92yp
t44ntqIwwKC8Jc156RgXNtv3ZAQ4V2ZPKh/hA6V8bcrFph0wIoHEAVT8tfzVylQm
R+oGm7LlMrEBYrxotQJCnF3aLOkeSbW8atjdF990ASyVCT+JzOk+cNT96DKncUQx
V8ES3F4CO3jlqgy5PJcLK+9oBPhkINsuk9RgQUTkKbj8Rgpv9YoSehkyMuUemREW
HiQOnLMBTk71b3ekY4EKXhO+/FHa7q9eQ3SF+RXehXXpaVK7Vx/8ig+aTLEGeepm
5Rxeg8g3hYOYGRLZd8fIzosVdrf0tG3KYxd/qL0eNZyv7ZYi1mi4a9W6lSjP8wNe
bbBva88tSUgOfEprYeK38K7/Ya8TOLFW1YBC3zf+3SU1Ul7elrEhsGDs6RGJPXQn
tHFGgVZP1+FoFmJWVzgwStZnLcAHWlmBnsqwbE0/jjSruRMgVOa/8Mbt7t+L4dLP
oNhV7kkFcrFb9YYA3sTGx3pa1R6oa60cpQFCl4Qg0uqI+QgwwezEvu2VKG0oVV/+
VS4m/qfrIHGcgd7dpb84wbdZmz+51y1sEFFjnLJzivE1wP2kPEySk2EOPzhd8vXi
NKug0xGEEdkylrPXdtgzLLs4QdmO4STh1DH3hlqzS4+wmBD7IM00j4bQW+gNx3MR
5IcEdMr65hOGei6V5WqYbtCzXPrgRselRWzmMj/z+4e7LEG8xFeN6vWC7LbzAFLF
eL3HFoGnwB2xqVnlHNJ2DHODXy6nVJxlkHgNAGPJIx2v29io0vfDI/xn/PUFrljT
hqk8Xj/q/Wpjgs5L2Wh1qSsiyXawTc1XODMjeQbCcbuaF5OYaFU4g0MOMQkbXmZB
QfTscdX+hj/8qMIf4o33CbeiIJTSCwjLEywiIiSP7tazsxhUykUI2heNptl7I1Af
A4T5HrEgrIRPU0dVzNSDLbll8ghdM/mRSBFyKKw6PnraRFi/CMsd+ICKNENBM7Gm
Eg6u7rT8x6QCspi6G9nskAuANTEDUI3xWM+5QVHEPgQmvSSMVhiKGYeh06iwAm4g
ofWjcsNdRLyUarDlreE/svB+MUYYitGjPiDOhcSip5xRBGngSG9L0fCKow++Y8Yw
mIVlf1J1th0XokZ0vkv1PjdJK4kDszDmpyxTaFWDX7BsN0IpARzxp7wsKCTgEVIZ
7fzxY9yK1BwKbN9RvzBaBNiSDZsH1DdhG94bBryfzLrgFuFX2xwHmqMzmth6jvyG
Ut94+0VeRf80C4xmndS6Sq9maYHjiaPhKZmIrcdbb7JQkeGdpOrfqqqgGzXQJJ7J
3NoO1Qwhl9abUe+BxMRb9HRBlVm6ax35/hHk1A7xIIQ9aJe8FUQdSnzY1cj8uOdo
KDCdp4vTSTTyJxSzkBoeQXXPCl+r4MdpmW+ZW694qqTVD8bZ5jeUJC0dB/vdXaoq
icUF6qpR0JXFycJ8to29Xa+Ph/Zw3ERNKAcOOt2LNtwuVp6mIBIzS/vBs+bU2hak
FFjrw7hz0q9vMZiugREPnh10QUQUFrA7gr1cGrLWRGURFvSBOHtfLky8EMhWSuuU
MF9ZhUg13APBf/v1z1FvO72QqN0ZKT7uHEG2vTIAm6SQYBFk23J3Ga3po/twjiJ5
x2Vzv4uMDNUdaCwwelzVh3eDcO9D4t4rBemvKJa3rk9gCEUK0D7t4ATtH3pFazdQ
E3PHibLES5NShqPD1BcR2lMfjZ2L+MoSrDuvlAyNk4gxrp+D7Lx+UxrBHnwfFWYC
du/Ryw3Nhu/Qqabn/42OKcgu10Ri4/U84IjVeS73i7aZTmdJKFTRdouqWmQ5lVpO
85xTf9yic0P8Y/Phd64qJtT/kV89AK3PgfeVi2K++raxuMQtf5KHehHS7z2daY8N
QbYrhzSltwaG/OYsydqgLeuUBaaBU/Z9Mf/ZGaP0sZ/x+zAL2rw+fMxGV3tc+DXE
BwO0M0p/qNW2P7NdY4NemFgoignxo39XUPT4+WnQHu4ff63XjWpXHu6xQwWSoioU
U9X7GR9tY2QrBE2x7CXpIRuY0tk3D53aSUY6Nda2B7CbdfaHzrFN6p9IEmNVC0eu
USruaiXCg7mCFuT2GmuakxiZZSZ59upM0og1qdgaIjc2Jt6yBZ/nn2+AOTH7lAce
rDoYM9x0WorJdbT0XEaRumNqgnOUlz7qiKujzI29qTKf6KNPqKPp8i+3FDUBMDFl
lc+goDAIsjL3KUR8PTV3QvwkgnwgUnzcznqfmYtI3VmdD7TDgZYPDkDweQBulpFg
8kJw/ugwLz5kWiHTeSLdYgmCwUNFkz0bo3j6L9pb5Y3DmkaIv6edKBi+n99f6OZg
lOL4w4ISxCsEeDl9O4WdFAyvadtNEe0AO/C6vC/VvhPyOfPYxfHhX/qkARPENk0j
lSLOPsLVFnuI0fhGrBDGKpDarIatznMIkXxuNg2B8VkMSGo3jWwraVWk86u7jyWa
KTs7pj55NEXUKfx5lvIbkrsxrj6p5+bKqsyCkx9S9Z5Ae0wc93VNMLOjmKFyFwbd
FRc1GJuPLUDEcKku2fINYD5PRsevOrsWuYV7jjq1vxtE/WHvfo2Dm5hAEZIT5CXz
TFdIjzq3ky+ADWupR3sJ/cDCC0rJDPZ0K6avXccLFoNAmx6yTiiJyOkK+b2bTf/2
xLBVFeFdgLsDu6uFfQgBxM/jwdiHxQlJO5nlTokxTG2rPvQQdjofZmukZ8t3YrlL
GtzL71iRicdOwD4ELjjGG989bBJBF0DADfWqswuPucwXpdyUQEsjsMvD++RosA4g
e289aZnD4UIKA5WiIAD6rnJF2ni+AlTODCca3q9dV5eN6N388yDlNGP6gqLTnz9d
SvgXKsRUWl05ie9rGdf9H0UHsdGSziPrGEj87IxGuYEP4IiwJQGPoGSQv7AzZ0WK
KIoJ1/CfIbC3sGkUXQbTCU7AsaSQxGStQh84j6HPS1T3KAnwQ637b0RS9BEQQKQ6
K/y9Uh7Yl9dNg1jczyH029w0+qy4AI6WNs5KMGwqW3mts4AGgiWMFbwn/+OtcLPP
lWNotL/3U0KRDbm7eo/KaWsEjE8gY6XRCYS/qKbmZBqaZLgkW2sWVpB6uxOq2bOT
/qoRuSOlv1xSczoeXPgp24m2t7dzI5+tEi/8HA4TaMoiJRtVbNPWtBZfee3brclJ
1tltyWxVRFSk9hU/arNFga1Hes6Or1xN49p0eyMok5aMUDAk/Lov0RVijv5/l0b0
tzNt6kLbiYMthLhoakY8oFT8I+H+JTspYuPxxyQ7T80ktIFmxgxzECx1eB3pFgiu
pGpmDOca/zSKhSZYU7Rciy4LYAxHPV4avi9oLnSDtzP1xAvXfN5vy+MuEO0eutrB
n0B6QJ9Pr95K9c8Q8rRpVgaIvMpK47fC6E1xdKA84tQGa6GCvDlxZrBTBZrKS8+h
L5PrVjZDMM1ByvBYiheW1VISUmutttyQoUSPvwSmtwhceZdQu0YaiH0SFqWF7hU+
eBlyVFiNOfLf9WN7gyptm4awveUq7ieo+f10G2P1czKYc0xuBIstBNIeoiCLn3rX
zy0PKv6RXcW2RqEossiOOJKML6StEC69fSePeFBt4KqW9o+V7x5gxkvkFFWRtMCE
TCLfeBdUs2GUB+O7kKjEb/X42oKrj1wHWi5b/qTdClsE+hoY/20LDuYSLGBXtHYk
ZiS7fLqDGCOJbYJlLGwnA4H9Ryb8KwwkbNb/gpha4NTtGo7lp2HY2EXo8Q9eVepP
3gspxdqYC0W6b66CU1esPVTBkhz5RPucEuv1wfrsA9YKRlIjVM0qs5HWcQq6vT4G
JF7tlpjgm3rvQhQGi2NUxckiJWA36HPBqJEn7OmwZEDlXusPvOAZXxU67KFwuDw7
vPkZ73af5LJZIbBDmK6ouiqn1W3YC1RzyujSzXnyyCtSdz6BPUrYzkgzIa4qMUAh
YKtchFx13BuyWeu15QT9BEXVfiuSdfoVUwnrHTcjM+XLsfj1DjAlo6K+aRIFIkrx
1Po4eUBOKdJQa+95vbaSwaxLjLKNTO1kXHme9fO3FP0ntGck2n7dH/Gt7nYy4eb8
Qte8ZuQDuTENNqNiXXQluXpp+/9nuHc3Y3LvONzSVpPYdnpsBmVIKSTsJEAzVudO
A+eYPuJ6UJt98sgalpP7++FDzcpF/OyLHfa47dXXZfUl4tne1FM6BDVXltcr5P2X
K8ndv2/oGj9o6CZSnnWK81BrZek1YBfQO73SCRRPlxZb19cZ/NcackaFeXAUQpjE
nqWM0WQELuFv4tvYMwev54zC/I6UWYnrXCKl4iqD16NBqXRpOrvk6PjWf2Cz6NgL
peV6d07TipJz1htJStCaoOmqzsZd1t0qlNVdka1k3tuJ+ql/VuiBk7w6B+KvGMj1
cW9ExXn1wzMu5fG8B+cxA/KvFFiY7dzGa0bWlh0DabGaxITUjyDuUn7yIkEqcqHW
oQmRpJMi+cwPIjE0mnxf1XBGIaT3iJ8iqCKIz9365g50oFsFyJrEPIfbujuNuKPi
6EvpSP88cTSltFU2Y2FrqkuI2+qHbJqNHpzYbkodFdfzwuLSV2alGuUCSTCibLF/
QALnxdEBkkADjL5hrWietR6tUArPZiLuYQLMeJtYrSbXz4iHTSSH7jYnJSVupO3l
68kaw4OCqWK/ORcqH7owkZY09R7PFQ9du1PgTwkMKyqYk+IGhIxMO3hUneofbBmh
uoiuSlNR/Gc0u6PZtickKMYWtnNkn2X7zUSKE1w6/jHkdrcQi+mk0GaEGSjnbjbX
AKVLk+rInM1w9+IozhJeRpuGd9hYPB3HpgV5FUzli7ih2SaoQuNjMjkwI/Y9EXhx
yPnoJ5Db3nvEhHRcsJFLdNprSpY8A+RpsSvCL3Q8iO15lmuTQDSsP6ScJX9IyGil
53+h6PirF48zqvZBYzPqObTcfEpk5RkHJHz4ekYXg6fc0sCqb5C8N13INWvkYM+W
3zp9thitfZpgcE5nAbzy/hs4fu7ux7QerXLLbd6akvbfo5ElgvCHmBKJlwaFo0/4
S9B9D3vOhCZRiYtb9QbeYKtVr0JgFiCT5d+NsneDGDmZ/oE7SQgebf0rWLeqiGr/
/klHkPAXeVZkAwnC4ch9jfpioXoDcrHJ8OQZ9jHAj/yan8alFC3y8VjmDgUPVZHS
B7UAVOak3Gd4tbO5Y/CR4y8ROvtLIrpFU/0vwy+q8ygZq5JWLXw+gPCBe2/2o18B
l/Pab2ZRRjHDDlWVJN9/F80Fp4gArLD9jaZ6RA6cuRa5b97v8SnEJeVTeTmX/AP4
yLSrpMs8fPOeTu94LW8Ta2gJVt8q4GdRIyAfLJY16v3ymWUqGc0InDVrt4PVQblF
Of4NsAT1tRtnDbmHae4YBcYNjsdWgQc2KdMUWP/Gn1HtrtbUfbWTLE5Lsl6F21Jv
Tw1j+EtBtCwt4iLplLvUMy9FJ/uMBQ//sVFjkizABtBKXS2D+NrRNiQtUqJ4Cr6m
9ypnSQqgdtmpIuWaYj9PVympuzXBDLMMDJVq+YtB3+ViTJIAywQOE8L7/qQKgg6D
+88AvYZE24Diwi4FHH0z1IS15C5aDWGPkS8flJM39hQdlyoiwmcM5laecqWmTyN8
wPU32do59irsDUl81ESOTXXKLJBWKM8I59JNVFJwfaMFb5kLMwGzU6i77tc7rurQ
N6aWme5Ve/8EavHhuinDFQIRiP+UIzLWUVex5WycEcG1Nj191hd1LLWJZ4Wf+0eM
6zdwr9/5pZp8qTi3SBUg8VCUJ3TJx5eCkfm1MvHm57ZGosKXkndL8XVxcz3s9ixw
FIXVc4RQ0cxkBZQsgmBYYceGXD+LtheIUOkdT8DGBCUtgBvzS/7YuUsg5sGqu+yH
JVzLEaYyA85wwlHHBgTK7tyF9cg3ez5bH8x6buSp7wQpz35l5b+fMwERn1bVClzk
M+6Is7E8dxrsNEm1P0rMBm6hepjX52E53dssuaoKzoRuZ0tmvqr443egjlRZbCup
uTTOU1IRJaIy5KLHkdwmuWF+r0Qr6tR0rnUyEiLm0rwwAjC2rVlN77PnfW/iMDRh
GsBkfn3ebFdYP0aMhae08f5FJq3f0jPehnVZk9qEeMFQUmBqWleAl4d8BwBMZcRb
Ci6e1eiLB514nLIrQJw8l7Gsxmpxl+Bjr6JAZ7AxxHCKI8F0sr1ncAed3GlptNma
XwJjZhpvCmrT8FUPtgVN2dK4IfXugTWWQ0T4B8YxYfdNJw/TXrTu3zkoEAcVQtM3
0+/1jQHuA/eT379oXGFrRdau+23m9xXVDwHW5LBdaBqTBtitr9ISu8ezGRTjCLEi
QZuNioUr/CeG55JbixsxSNrT/FEM2eVfd3GSBANIRGeYH1vGa57qMtB2FG1gQ4d3
Oc4ykEDy6Vrdni2m625/nIDpZMe3So5QxiO0tE8+4vjahUtA//1teJB3F/Fq7K0v
i2sVgElqCyLcbgLoPWFKsbnXmPzRs2sO30S/8ycNJhwlfCMlA4VYWKYOo2IdveXt
7hrDtkmIMfCfQkvBD94JvNtFwEGU744Uy3nIq1BgbSofBK3FJAmparI1UHGlGPGA
fWUq4sFN2rbVEkvH8xicZ2cnYY4NbgRyvlRvVybMLSNb++Ux9KrRUetX33MdDdwI
eaye60GkS1FdsqKUtl8rt6j+5lYL0zYaBQ9IO4SDH6Jkp27lPLvAuix6C7258jx1
0hyyk7M0wQH7my5lb86FgyZLtfXzjWpR8bxyx5qBYKoWqOlyY7SwK4lqDHHHt1Jc
ZSYLiUqrsd62BMeuCtDn5ud8i0Ycrhkk/uC1ABrVW5VxUtXtAhWdsEdb6+qMDmsj
aGxYOKGt/51k1PRf3VVBRjuOsw1Ps8C4Koi72zrA7OsHZGyGcWqlXPdX+WcIFKYz
/HI2NWtnt+ytPzOXR3JBJL+Gdighw0fYuLFufZq5s9aH2lnY6pGQ+oOJqZCKKScX
G5Nkjwvde0svLrIq681T3jZ+VNnlpYwuZoOk9Xw5ccvJ1R6IRwW9OJZz32+db8U5
vq63ofebtWyDI8YKCkHriEm5Wh6MiFdxadnaXLx9lS96Mq5FhGkTopiLqg+bdnZd
aGa5YGFCjUqZwvtlpczMIkeNKaUTV+X/arbBMHE11oFN9yGNlxgjnHOfg5cC92N8
RK0Kh1TIA3FcToRI6+Es6kc6Zm3X5fQ7JIxfbuO4pxXS2xB8O1LIdh3wUQsaPLh3
N9Z5x/4xy36vpBFlbDbSKj0dohXb6jt2Rvgx+U6VfgXfOBA1Qwk3LOR+nA3kq4KO
W2gvtVterGpovnGVc7+H12k6xXgyqGjZNDbHFFl6zZ9RQnDslspN5AZb0vvcc7pt
3/mESeDehBqXsL4Ufs2Tj0RCTwzA8ih5dey3zsEL0pMkXWXJdzFltsMNTRtaZTsw
jjcCbByyO+lUxARD+hAVBafsCOe3v1JSuDnJkdeiF3AgHAvZEQWeTd/M+978HO9r
fIh5mOnV9NG2PQb07QzaEOFGimVwQ2tFUQnOJrYobVpi5snCJ2KxBvpMZqrM4VRR
wYBVV8zqN0UTpUS8z5e3UM4eDLRM+WfhD6yViMxrEiYZ+xd95joueTnCGCc1TvEv
Iyk2eRyV8yAWvQUfPBrpnkvlB0itZB666FCXk5pRlyxa8JMsmiUcld4NnYrTTUvl
kzW/8OquAAHE5JXRAl2VQvBbt2hq+VSBNgW73aZ7WQsFSIzQW0GnJekhNxZncp/B
FevBJvUO+8hoo422+OLQZp/u8VTxC8jqJMt9zwVz5wwzc3qpz5M+WA3wcAtUb3gc
HtyIl3yYd5nGK8doQg5RLnCXfVdlmotmyRMJuAG3tbVgxzqqpolFMwTUdGIx51n3
S/RHGliZLax5yyLPeln7S2HIQHzfgJiZDKajGmFxTuAg4rO4sBy51HBftEUQFYvW
yDaBgrc9kY+8SGsgaUZDRejok7ilFe9RHvqwQszPeVcZ2Uf8YvLmRZ+6NOVHtKyK
+aFS5onvE1zuXApHazz8gA14RvL6VGSj3uooAX3xgKL/OKoqtqYELqgnkeZubqK3
Nlji8emHsHUs7xsKr23c2i3MuzUX/z9d0bwO7P1htPurBU/bpEKO06u/bEjmPs4p
UIXnC2GItbizPgaCxiakUYRVRUY1a1pe0rdTnK1Ne2qpthKLMoEZfRmeEBtxHLy1
uAAoucJl214OIeeM9A/dSj7GyZjeYTi4Mwozy9PyKWFKkohMrgg2tgAkqfYHrBEB
BQB03mwODmWtcRBw3WGLE2+OnDr/d94J77DPFrBT+EwiFR4aR2eyKQtWHTUt1BIF
1xods4N9K6/lIgVX7c5xsagTTsLyh06ovtngB60KfkyzKOs75gBT14Nw4qZThZem
dVUaxqYS1SGxD0wGD8Ka7XHttiKtlBPkliGT8SbtAw9gxeX0yK7ZaEctt21Ka4oC
1TFv3lCWx1NNcWxTclWMwNvCaXXuOkEg1FTmVUFrjP+mARB9T4WcBmvMB9VvrarJ
YMy9L8ltEGM048SlexelPFgeZ+KADiv+YggS521gSxCnOWvmiAAW1pNE9LgfaLZ6
Q+gz1isWy2d32OS5/b3uPcBT+yw4RBiFPCw7/WNtghKC3kQ1Nu6SkhRCegHblrwN
YOv/g5Wo29Q9hsbC6CxqRKM5RZX7QzCOU2fkxfD43gIsnQTSzeFY0jF9ghyAsPYs
0xBsa387hyd9brY6KDFCuWutq/9rZIJtCNIKKNH4ArGYkqRicjZGnG13TBANAuoH
HhuhCnfMYjK2jtYEXs1qZsaVEci0MFPkuyqj5PCXTYg8+TUiI3716cbXenSOGR2N
t1DHxPHi3skOUXxCQZkKW+bIWfxENEwMKm5UTO3bRKJiNCVLo3+XomUe2lKr+ep0
/RzHkk/rHQLvmPfxcknZpgOEaCOE49oAZW3HuxuzmhPnpdD8w/1aovqxYJomlvi9
qM8Xwka33qNjol4oy92F+aQYRoVM6/Tu6GK2+5EzKBKnX9H3Z5XXKT26R5evq+3Z
849O+h9H6ABG8J/Ya+FfuiFToxNOGDAfJv3Hv/a0DS5DOBULy2KlO1hNeyqvWmwS
tzElNAIXy359UT8q34RcDzcYBmMhCOAhkFT4pGfnaoARKzDEJ3CAWZ/CZtNgjjvT
TJ/n+k/7Vsu3hv3z41tsFj+fgzWbUmSqiCfbJ81e7RgjQZNlmLQksJ22kQZBzd4y
Ymv47UWe7i4ZCjLBds/eO1WjZm275PyVPqPFCySnkUdrlIlCDz2SoLOEmXus/8py
x8JrkIyvOlD1r/eTLpZusSPp3MQgNCVSnQoQXfGbqteCNZhEhcCOI9BTow1UG2pN
ZV/8D6tuTeQYTLO1G4tjhKXvG3dubltT2ejT4CSy1IRZZM3JCgnsGyGbq/Y6FFdh
x6pD+QociqtJPHArhKFrUyr5+/0WipdN4R+8loACl6DfTQkNRHN+qWg/K9zv59sL
1b/5g+8TOsA1Hj3qGheYEgJ9hd9T7yRmTT49KsDsocT0L4AF8ZbURkvEujy6tkjg
WzJ+sSdhxAyn9Xqft+vTo/XKkf0lr5fqPAUBCJ1C26M/6SROaiOslRbgAdrz9DQY
HAg71SBJd47JQPBpp+5DEgZfyJhIC0Fa9OlN2ENOefymPAYCNIAqBBXwIsyMDlSb
A/Lg7SpxLY6UZemp6HW/b98CQpvM9X9ozP4FSFsojpg4e8S9j1CO9zz+ZqKDx/XC
FunhduJdQdD3qgwe81XpvlmVQxwDRZ9YjNTVxBRpQwKtsfRx/mWZyimsHm0pHZzb
pWVvabdLz0UnhuY462tMmWdKybSrA2i0UdBvuUHid9uN7/rimpO5Aec3kGhYDkDO
q+scIe38eI48zxMyeWCf+B1WHk1tX2wnTm3ixyifUp+vOB96rbTnfq2htbyRxV0V
oGeEippHwHzJK2hGJGIBdkmSbY4NYobFJ5b27nRGZOczctFI94XIOV9ZQKFfIKo+
IjTFHPu+UKpcl7nFaD2TFsI18scYkPpwWnObpOBKdk+xNnFzYozCdGkWePW9D4ug
FzmmDK6+W9xt4DBUVNzYwVt1pdVWA5vCcfGO8XIx2risSUQbHjYNNguidaKNyfLv
jLJQay4u1bjjz91CBDX3vGQNl9hZHdels2LvQyDjti/cT+WzbDyVOfowHMvmHYFm
jTTOPC5jPeVZrYh39nwnQaBOEY4qkkTkoYqVZoVTOQwnBPqF0M1GvocTdm7gBwYv
1RSmiErz5uZdw7V0zdvL5bZD1yJa/4BxTFwWCCNgKQxmyeiIeyejLECifF2xXavb
mnDAUbF/QaW5uXx7Z7NPfZMLKfQ+rUItxfyH6uj30hjZPZsURQveBytyZ2Rk6ePO
AO6Y1FSggBpWKpyKFQfK4f+Gg7jX9q/4GGTnDnTvqNNbV+dyNm0QWfmHLqejvB0i
WeclwYURkEjftZ+/F+rd7Y+kZeRVI+yzZ2KG7WStd1oZ6Nz8+965U6TCRRIL/LmS
3984nrpI4WKmgDaMM1YaklIi90RfOReN5HCfRfblRY4BmMWqgjAG9S12vkkm1FvG
anLYeRR3hq3J6BADBvrfeu5dGzjkNol6LfnX9QsgAdvE83NdTK/VCyUUbhnYhlbH
9Yuwj/TIk+wA6zPAVEbeG0Evn6HCrruzXg1pwoU6+TMPYkZ7tXaNabDYoHCVZCxb
xlcS9MG72RXNBjLQMii90aQeItsruQWQiVlQVPeYF8X6AsZmJ3lbCzYlT0TY5mZG
2sjvutHRas6R4qXw36WSR4cSM5rys4Fctp5WjPIBaRRHLJO+oblHO+bk1C6btGsZ
Ge5MxOyRTkQUJBgzLrn9GGbnyZ+Mh9B8NyM/JRnSIK7HznPZGRx9JGrLSBgv6GCc
RyZZdnz03VijyRhqaVQaEgne0Dw5yzZDYJdHpRjh79Iq48I7F4M2IovlqJjpCZRC
9YtFUWXapiGma6vChwXl0M/D6oKWNzPMCKOUUTfhaEFi3VkTlt6ct7+VFQbOeWaA
Ve1FBs/KznRLnAh7AVTJYFYbJ/MaEzLhkCkaakhctmvxZ+Pbmjwvlzu3Oe7FLxmm
1eSQCMh4QF8IKEdD0PzSCvTnJlb64K/4LV+c0kp9JSm4s6/n5gSCvsUW7Fp+n9Jv
34cVGvM1wdgjGsMGICMA0SjlkrKfKZ3zOKRFdJvnluyfBLJXzLLd8z4D3NLCgRit
3rg2MpCsgol4p5rPb+v8RhaxL/uFG1R9N32oBF6ApeBynmxWT5KDROLhsZhvvN6S
/2qck5115aMwXL297PdQBZvbn9Kae5St5myt5cgSu0S55pChNc1bA/aXsUEW9jgS
TCBGL+ZnshEqKO3JkIXWwebG7LG4SAlyaQyqlWtDnmTU9FUUqV6GcjYOjHZcDy+x
n9nNZHgz9922XMZvqv5Vu4/cu0ocf8+PcZy3W6gNNsewxZ4FX2Tz+raZs08yvyhU
4fQHBbXHlffbL/3QaaWQccWoInvxpsIegyMR9Qy2Ne0vDeKQP2FrSVGk7KDlgsHh
J8fPSAjjYNkgtwVUmpoWkzusWrb0xRIvYkyDNmJPGwFrykypBavoS56fSSrAzvBf
hkpWSOwxovF9N+BTH3FG8g5x6cTwGnbyNb7yvM0Ywi/A6KATaIQl53JpozckHLM1
PlJd/sQV1WGrx5W/6djl4MjEk6iqWxvDa5u5UYAhBFFfYxIW1GsB1t862UqJopU4
MPww5GclM+EEVHVAWQAQrIqlLQHfb7dXfg3cSWQ80KuLxixoX4gdnHu0mdA04Odr
/lp4DT0U4wErFgbBqY8JwSwXBfMN70gnxlGgm9/fvopVFhJq4pIcq2ddnntdXWkm
L1nE/D0ubTrmJW1DYGqft/uEdEwgLMobPnjZsnVFYSXeeW6i+UxVK32li4SXfJ2+
Kbf+4kJ527S1USB+43eG+vjZRQnA5iMQhFOM4YaJ0WEs1i1kudeSEObKi3fmy80b
KNECR8qJK2MeId/DnQByFDwIpf4wHxQPi7S0IkwJrae6yO22dmJNrFmz0CQ3geqK
wbfJ9TmRxAM+M7A3G8glQ056EVFucXoyJ6aT5f7q8uKqDOOamTxF8eHBKZcPD9Am
TKg9jHXtYINr4fhZnzpRTYM+2Xifpqv72ykJP9ySHaeX9bQ4oPzyC+YJknDjHBxX
mZIVx5rpKXvJDVU4+0nARfvG0c8Sv+UTAzjaA3r7XfFxCNoj5WQZxp0TuhfeKu03
RPnWRpZmJ5nCI5Oz3JiK8mXIoZ2VsrSoZJx4kJLjnSEYv5Hx2/I3oPBxC/vVYSvW
jUVXHaGeMuiA2zT8G6SWX/wciIdzCwrDIiAY2H9jtD8SejmNlCPloYIXruje8dTg
Y9estEa3/ocI/IB550xfM/5NRks/3Ip1a+/kY+e7zNBqZQVAoLnf95Z0fmcNEcZ+
eQXNMV4Lsca0OHmjB8B9NZBil04BlfrmkzE6MjHYk6wPTS3ph0BnyYupJcsBFuoL
fDWcahN9Ne35I6BZlXp1tmCbtaeIHrOMsK0wJNRc7DSHZ2+c12bAdWP+gaT8pC3e
AgFLerani5AKXl1Y4DsYwThNmixTOndJ1TafB2NhTAPYzjVeoIa96RTMDipWmlh8
qn6zxKKdBmvlsNt8kbCvRjDBZpiHhu59/qRhuuSOBUk0s80djNqwJAzEkx26p0ux
gdRBr2ndBOUl2dms9xAnUnZ3A9v/gzxANc/gFzrzbHQObMcZi+zmQus9idcDpeTF
1ayxxEhV/OV746TE8at2oKs0r32kmIukgZyGZAjcgPmRbdoYoI0OdOY7fMyD1TRu
nVAE95s7xIJP8/meMSHynlM15mYfVW6r5EjtN5HOv9jRln79rKB3SsEbTgxzmInJ
l6Jan72iT7WzY/FrIyQh9/k8Z7m+KZcNPAP9Uw1MqVuXFmJ2Pk5Kum3ARujdRSoy
aJPz/QyRMHt5puvwsXY6h8SQYYKQRSMoMoZbQjkMnnpGeNfUaQILILXzMbpDTXsr
fJU5Fdc/x9ZPiVHCJxIgO6zXF7ZK9xtaNZu1vOEk1YyIUygAQxVbeldMZBCZ9sz+
zIo/qLjud/eLKYAGuwgGpWVuLhTujAdIf0/8TMr9PbLNBJoLHWxGrlszeSlJd2mU
DbNNvRUopXMN9jnwvh9IX4mVVLNCZtUnuH8BNdowMF5+GEaEUjL9ZQF3Skfb27PF
MccFMBtXKux8Xi2TU/XcKAskS9jjpdN76BNCvKnOpwc80GEqxoOQI9UNPMTWEFmC
T0t2bc67BqmB9SHEyTndlIZlKm7VbugX0Gw+RmKjTwHZQ+ThA66nCNmUfmy7yrYG
dzj3wgGZPJuSHSk8wAJ+LVrJv3kpUEqGjRAXTIffTO0nQQihkZmPEBeePG9Buv3R
E+9KXeJdR4ork2t4JGDKtgcjTnGaiujrN/3+XbeufRC2QfyBS9tXS/AO5XA9SUp5
X996yE5KF8Qy+TTvxO1rww==
`pragma protect end_protected
